module ROM(
    input clk,
    input[12:0] addr,
    output signed[7:0] out
);

reg signed[7:0] m_out;

always@(posedge clk)
    case(addr)
        13'd0: m_out<=8'b11100100;
        13'd1: m_out<=8'b11110000;
        13'd2: m_out<=8'b01000110;
        13'd3: m_out<=8'b11101101;
        13'd4: m_out<=8'b00100000;
        13'd5: m_out<=8'b11101110;
        13'd6: m_out<=8'b11100111;
        13'd7: m_out<=8'b00011000;
        13'd8: m_out<=8'b11011001;
        13'd9: m_out<=8'b00001111;
        13'd10: m_out<=8'b11110011;
        13'd11: m_out<=8'b00010010;
        13'd12: m_out<=8'b00001111;
        13'd13: m_out<=8'b11111010;
        13'd14: m_out<=8'b00001111;
        13'd15: m_out<=8'b00011000;
        13'd16: m_out<=8'b00010111;
        13'd17: m_out<=8'b11111101;
        13'd18: m_out<=8'b00001111;
        13'd19: m_out<=8'b11110001;
        13'd20: m_out<=8'b00000010;
        13'd21: m_out<=8'b11110110;
        13'd22: m_out<=8'b11111011;
        13'd23: m_out<=8'b11010010;
        13'd24: m_out<=8'b00000101;
        13'd25: m_out<=8'b11101001;
        13'd26: m_out<=8'b00000000;
        13'd27: m_out<=8'b00001111;
        13'd28: m_out<=8'b00000010;
        13'd29: m_out<=8'b00000110;
        13'd30: m_out<=8'b00111000;
        13'd31: m_out<=8'b00000010;
        13'd32: m_out<=8'b11111100;
        13'd33: m_out<=8'b11010111;
        13'd34: m_out<=8'b00000001;
        13'd35: m_out<=8'b11111010;
        13'd36: m_out<=8'b11110000;
        13'd37: m_out<=8'b00011011;
        13'd38: m_out<=8'b11110101;
        13'd39: m_out<=8'b00001111;
        13'd40: m_out<=8'b00100000;
        13'd41: m_out<=8'b00011110;
        13'd42: m_out<=8'b11111110;
        13'd43: m_out<=8'b00001000;
        13'd44: m_out<=8'b00011010;
        13'd45: m_out<=8'b11000100;
        13'd46: m_out<=8'b11001000;
        13'd47: m_out<=8'b11110011;
        13'd48: m_out<=8'b10111111;
        13'd49: m_out<=8'b11101010;
        13'd50: m_out<=8'b00101101;
        13'd51: m_out<=8'b11101000;
        13'd52: m_out<=8'b11110110;
        13'd53: m_out<=8'b00010100;
        13'd54: m_out<=8'b00001010;
        13'd55: m_out<=8'b11111111;
        13'd56: m_out<=8'b00001000;
        13'd57: m_out<=8'b11100110;
        13'd58: m_out<=8'b11111010;
        13'd59: m_out<=8'b00000001;
        13'd60: m_out<=8'b00101011;
        13'd61: m_out<=8'b11000010;
        13'd62: m_out<=8'b00000010;
        13'd63: m_out<=8'b11101011;
        13'd64: m_out<=8'b00011100;
        13'd65: m_out<=8'b00100101;
        13'd66: m_out<=8'b11011111;
        13'd67: m_out<=8'b00000111;
        13'd68: m_out<=8'b00000001;
        13'd69: m_out<=8'b11101110;
        13'd70: m_out<=8'b11010111;
        13'd71: m_out<=8'b00001111;
        13'd72: m_out<=8'b11110000;
        13'd73: m_out<=8'b00010001;
        13'd74: m_out<=8'b00100101;
        13'd75: m_out<=8'b11101011;
        13'd76: m_out<=8'b00011110;
        13'd77: m_out<=8'b11111101;
        13'd78: m_out<=8'b11100110;
        13'd79: m_out<=8'b11101111;
        13'd80: m_out<=8'b00010000;
        13'd81: m_out<=8'b00101010;
        13'd82: m_out<=8'b00010100;
        13'd83: m_out<=8'b11101100;
        13'd84: m_out<=8'b00000100;
        13'd85: m_out<=8'b00100001;
        13'd86: m_out<=8'b00011111;
        13'd87: m_out<=8'b11111001;
        13'd88: m_out<=8'b11011111;
        13'd89: m_out<=8'b00000001;
        13'd90: m_out<=8'b11110111;
        13'd91: m_out<=8'b00000110;
        13'd92: m_out<=8'b00000111;
        13'd93: m_out<=8'b11010011;
        13'd94: m_out<=8'b11101110;
        13'd95: m_out<=8'b11100111;
        13'd96: m_out<=8'b00100000;
        13'd97: m_out<=8'b00000011;
        13'd98: m_out<=8'b11101111;
        13'd99: m_out<=8'b11101001;
        13'd100: m_out<=8'b00000010;
        13'd101: m_out<=8'b00000000;
        13'd102: m_out<=8'b00010001;
        13'd103: m_out<=8'b00011101;
        13'd104: m_out<=8'b00101010;
        13'd105: m_out<=8'b00101011;
        13'd106: m_out<=8'b11100110;
        13'd107: m_out<=8'b11110001;
        13'd108: m_out<=8'b00100101;
        13'd109: m_out<=8'b00000011;
        13'd110: m_out<=8'b11011111;
        13'd111: m_out<=8'b11101111;
        13'd112: m_out<=8'b11111000;
        13'd113: m_out<=8'b00000101;
        13'd114: m_out<=8'b11110100;
        13'd115: m_out<=8'b11101000;
        13'd116: m_out<=8'b11011111;
        13'd117: m_out<=8'b00000011;
        13'd118: m_out<=8'b11100100;
        13'd119: m_out<=8'b00000010;
        13'd120: m_out<=8'b00000011;
        13'd121: m_out<=8'b11111100;
        13'd122: m_out<=8'b11001110;
        13'd123: m_out<=8'b11100111;
        13'd124: m_out<=8'b00101010;
        13'd125: m_out<=8'b11111001;
        13'd126: m_out<=8'b11100110;
        13'd127: m_out<=8'b11110111;
        13'd128: m_out<=8'b11100011;
        13'd129: m_out<=8'b00010000;
        13'd130: m_out<=8'b00100011;
        13'd131: m_out<=8'b00010001;
        13'd132: m_out<=8'b11111110;
        13'd133: m_out<=8'b11011100;
        13'd134: m_out<=8'b00000111;
        13'd135: m_out<=8'b00000001;
        13'd136: m_out<=8'b00001111;
        13'd137: m_out<=8'b00010000;
        13'd138: m_out<=8'b11111100;
        13'd139: m_out<=8'b00111000;
        13'd140: m_out<=8'b11101010;
        13'd141: m_out<=8'b00101110;
        13'd142: m_out<=8'b11101101;
        13'd143: m_out<=8'b00101000;
        13'd144: m_out<=8'b00000100;
        13'd145: m_out<=8'b11110110;
        13'd146: m_out<=8'b11111110;
        13'd147: m_out<=8'b00011110;
        13'd148: m_out<=8'b11111110;
        13'd149: m_out<=8'b11110010;
        13'd150: m_out<=8'b00011100;
        13'd151: m_out<=8'b00001100;
        13'd152: m_out<=8'b11101010;
        13'd153: m_out<=8'b00010111;
        13'd154: m_out<=8'b00101010;
        13'd155: m_out<=8'b00010101;
        13'd156: m_out<=8'b11111100;
        13'd157: m_out<=8'b11110111;
        13'd158: m_out<=8'b00010100;
        13'd159: m_out<=8'b11110110;
        13'd160: m_out<=8'b00010000;
        13'd161: m_out<=8'b00010010;
        13'd162: m_out<=8'b11111000;
        13'd163: m_out<=8'b00101010;
        13'd164: m_out<=8'b11110011;
        13'd165: m_out<=8'b11011011;
        13'd166: m_out<=8'b00001011;
        13'd167: m_out<=8'b00001110;
        13'd168: m_out<=8'b00011010;
        13'd169: m_out<=8'b00011101;
        13'd170: m_out<=8'b00000011;
        13'd171: m_out<=8'b00011111;
        13'd172: m_out<=8'b11101010;
        13'd173: m_out<=8'b11100010;
        13'd174: m_out<=8'b00001000;
        13'd175: m_out<=8'b00000001;
        13'd176: m_out<=8'b00100001;
        13'd177: m_out<=8'b00100111;
        13'd178: m_out<=8'b11110111;
        13'd179: m_out<=8'b00001001;
        13'd180: m_out<=8'b11011110;
        13'd181: m_out<=8'b11100011;
        13'd182: m_out<=8'b11101011;
        13'd183: m_out<=8'b00010110;
        13'd184: m_out<=8'b11010100;
        13'd185: m_out<=8'b00011000;
        13'd186: m_out<=8'b11110001;
        13'd187: m_out<=8'b00110110;
        13'd188: m_out<=8'b11101011;
        13'd189: m_out<=8'b11111101;
        13'd190: m_out<=8'b00011000;
        13'd191: m_out<=8'b11110011;
        13'd192: m_out<=8'b11101110;
        13'd193: m_out<=8'b11100010;
        13'd194: m_out<=8'b00000001;
        13'd195: m_out<=8'b11101101;
        13'd196: m_out<=8'b11101000;
        13'd197: m_out<=8'b11101010;
        13'd198: m_out<=8'b00000010;
        13'd199: m_out<=8'b00001001;
        13'd200: m_out<=8'b11010101;
        13'd201: m_out<=8'b11110100;
        13'd202: m_out<=8'b00001101;
        13'd203: m_out<=8'b11100111;
        13'd204: m_out<=8'b00010100;
        13'd205: m_out<=8'b11000100;
        13'd206: m_out<=8'b00001100;
        13'd207: m_out<=8'b00001001;
        13'd208: m_out<=8'b11000110;
        13'd209: m_out<=8'b00001010;
        13'd210: m_out<=8'b00000110;
        13'd211: m_out<=8'b11101111;
        13'd212: m_out<=8'b11101001;
        13'd213: m_out<=8'b11011011;
        13'd214: m_out<=8'b11000110;
        13'd215: m_out<=8'b00011101;
        13'd216: m_out<=8'b00100001;
        13'd217: m_out<=8'b11100000;
        13'd218: m_out<=8'b11011010;
        13'd219: m_out<=8'b11101100;
        13'd220: m_out<=8'b00000100;
        13'd221: m_out<=8'b11101001;
        13'd222: m_out<=8'b00000010;
        13'd223: m_out<=8'b00101110;
        13'd224: m_out<=8'b00101001;
        13'd225: m_out<=8'b00001001;
        13'd226: m_out<=8'b11110001;
        13'd227: m_out<=8'b11100010;
        13'd228: m_out<=8'b00100010;
        13'd229: m_out<=8'b11111101;
        13'd230: m_out<=8'b00100100;
        13'd231: m_out<=8'b00001011;
        13'd232: m_out<=8'b00000011;
        13'd233: m_out<=8'b11111101;
        13'd234: m_out<=8'b11111000;
        13'd235: m_out<=8'b11110001;
        13'd236: m_out<=8'b00000011;
        13'd237: m_out<=8'b00001000;
        13'd238: m_out<=8'b11010000;
        13'd239: m_out<=8'b00010001;
        13'd240: m_out<=8'b00000100;
        13'd241: m_out<=8'b01100001;
        13'd242: m_out<=8'b11101000;
        13'd243: m_out<=8'b00010010;
        13'd244: m_out<=8'b00101101;
        13'd245: m_out<=8'b11100110;
        13'd246: m_out<=8'b10111101;
        13'd247: m_out<=8'b00000101;
        13'd248: m_out<=8'b00001011;
        13'd249: m_out<=8'b11110011;
        13'd250: m_out<=8'b00010001;
        13'd251: m_out<=8'b11100111;
        13'd252: m_out<=8'b00001011;
        13'd253: m_out<=8'b00000000;
        13'd254: m_out<=8'b11111011;
        13'd255: m_out<=8'b11101101;
        13'd256: m_out<=8'b11001011;
        13'd257: m_out<=8'b00010111;
        13'd258: m_out<=8'b00001000;
        13'd259: m_out<=8'b11101011;
        13'd260: m_out<=8'b11111111;
        13'd261: m_out<=8'b11011000;
        13'd262: m_out<=8'b00001100;
        13'd263: m_out<=8'b11100000;
        13'd264: m_out<=8'b11010110;
        13'd265: m_out<=8'b10111110;
        13'd266: m_out<=8'b11101100;
        13'd267: m_out<=8'b11101001;
        13'd268: m_out<=8'b00000011;
        13'd269: m_out<=8'b00111011;
        13'd270: m_out<=8'b00011100;
        13'd271: m_out<=8'b11110001;
        13'd272: m_out<=8'b00001001;
        13'd273: m_out<=8'b00100011;
        13'd274: m_out<=8'b11100110;
        13'd275: m_out<=8'b11001101;
        13'd276: m_out<=8'b00000110;
        13'd277: m_out<=8'b11010010;
        13'd278: m_out<=8'b00000011;
        13'd279: m_out<=8'b00001111;
        13'd280: m_out<=8'b11111000;
        13'd281: m_out<=8'b11100110;
        13'd282: m_out<=8'b11011111;
        13'd283: m_out<=8'b00001110;
        13'd284: m_out<=8'b11100001;
        13'd285: m_out<=8'b11100000;
        13'd286: m_out<=8'b00001100;
        13'd287: m_out<=8'b11011001;
        13'd288: m_out<=8'b11101101;
        13'd289: m_out<=8'b11110111;
        13'd290: m_out<=8'b00100001;
        13'd291: m_out<=8'b11011010;
        13'd292: m_out<=8'b11101101;
        13'd293: m_out<=8'b00011000;
        13'd294: m_out<=8'b11111111;
        13'd295: m_out<=8'b00011000;
        13'd296: m_out<=8'b11101011;
        13'd297: m_out<=8'b00000111;
        13'd298: m_out<=8'b00111001;
        13'd299: m_out<=8'b00010000;
        13'd300: m_out<=8'b00010111;
        13'd301: m_out<=8'b00000010;
        13'd302: m_out<=8'b11101100;
        13'd303: m_out<=8'b11101010;
        13'd304: m_out<=8'b00001001;
        13'd305: m_out<=8'b11110000;
        13'd306: m_out<=8'b11111001;
        13'd307: m_out<=8'b11101000;
        13'd308: m_out<=8'b00000111;
        13'd309: m_out<=8'b00010110;
        13'd310: m_out<=8'b11101011;
        13'd311: m_out<=8'b00001011;
        13'd312: m_out<=8'b00100011;
        13'd313: m_out<=8'b11100101;
        13'd314: m_out<=8'b11101011;
        13'd315: m_out<=8'b00000100;
        13'd316: m_out<=8'b00001111;
        13'd317: m_out<=8'b11111100;
        13'd318: m_out<=8'b11100110;
        13'd319: m_out<=8'b11101010;
        13'd320: m_out<=8'b00101011;
        13'd321: m_out<=8'b11111110;
        13'd322: m_out<=8'b00000001;
        13'd323: m_out<=8'b00001111;
        13'd324: m_out<=8'b00000100;
        13'd325: m_out<=8'b11010101;
        13'd326: m_out<=8'b11111010;
        13'd327: m_out<=8'b11110001;
        13'd328: m_out<=8'b00001000;
        13'd329: m_out<=8'b11111111;
        13'd330: m_out<=8'b11101010;
        13'd331: m_out<=8'b00001111;
        13'd332: m_out<=8'b00001101;
        13'd333: m_out<=8'b11100110;
        13'd334: m_out<=8'b00010100;
        13'd335: m_out<=8'b00100100;
        13'd336: m_out<=8'b11101100;
        13'd337: m_out<=8'b00010100;
        13'd338: m_out<=8'b10111111;
        13'd339: m_out<=8'b11110001;
        13'd340: m_out<=8'b11101011;
        13'd341: m_out<=8'b00101111;
        13'd342: m_out<=8'b00001110;
        13'd343: m_out<=8'b00000001;
        13'd344: m_out<=8'b11111000;
        13'd345: m_out<=8'b11111101;
        13'd346: m_out<=8'b11111001;
        13'd347: m_out<=8'b11101111;
        13'd348: m_out<=8'b00101011;
        13'd349: m_out<=8'b00000101;
        13'd350: m_out<=8'b00100010;
        13'd351: m_out<=8'b00000110;
        13'd352: m_out<=8'b11111110;
        13'd353: m_out<=8'b11110100;
        13'd354: m_out<=8'b00001100;
        13'd355: m_out<=8'b00100100;
        13'd356: m_out<=8'b00010011;
        13'd357: m_out<=8'b00101000;
        13'd358: m_out<=8'b00110011;
        13'd359: m_out<=8'b00011010;
        13'd360: m_out<=8'b11100110;
        13'd361: m_out<=8'b11110000;
        13'd362: m_out<=8'b11110000;
        13'd363: m_out<=8'b11110110;
        13'd364: m_out<=8'b00011101;
        13'd365: m_out<=8'b00001000;
        13'd366: m_out<=8'b11110101;
        13'd367: m_out<=8'b11101111;
        13'd368: m_out<=8'b11110111;
        13'd369: m_out<=8'b00100111;
        13'd370: m_out<=8'b00000111;
        13'd371: m_out<=8'b00000010;
        13'd372: m_out<=8'b00001111;
        13'd373: m_out<=8'b00111011;
        13'd374: m_out<=8'b00011111;
        13'd375: m_out<=8'b00010100;
        13'd376: m_out<=8'b00010110;
        13'd377: m_out<=8'b11111100;
        13'd378: m_out<=8'b11110001;
        13'd379: m_out<=8'b11111000;
        13'd380: m_out<=8'b00001010;
        13'd381: m_out<=8'b11111000;
        13'd382: m_out<=8'b11001100;
        13'd383: m_out<=8'b00010001;
        13'd384: m_out<=8'b00110101;
        13'd385: m_out<=8'b00000000;
        13'd386: m_out<=8'b00010000;
        13'd387: m_out<=8'b00001000;
        13'd388: m_out<=8'b00001111;
        13'd389: m_out<=8'b11011110;
        13'd390: m_out<=8'b00001101;
        13'd391: m_out<=8'b11110010;
        13'd392: m_out<=8'b11111101;
        13'd393: m_out<=8'b11100111;
        13'd394: m_out<=8'b00001111;
        13'd395: m_out<=8'b11100001;
        13'd396: m_out<=8'b00001001;
        13'd397: m_out<=8'b11110101;
        13'd398: m_out<=8'b00001110;
        13'd399: m_out<=8'b00010001;
        13'd400: m_out<=8'b11100110;
        13'd401: m_out<=8'b00011001;
        13'd402: m_out<=8'b11100011;
        13'd403: m_out<=8'b11110101;
        13'd404: m_out<=8'b00010111;
        13'd405: m_out<=8'b11010010;
        13'd406: m_out<=8'b00100101;
        13'd407: m_out<=8'b00000010;
        13'd408: m_out<=8'b00011100;
        13'd409: m_out<=8'b11111111;
        13'd410: m_out<=8'b11010011;
        13'd411: m_out<=8'b00010010;
        13'd412: m_out<=8'b00100000;
        13'd413: m_out<=8'b11100000;
        13'd414: m_out<=8'b11101110;
        13'd415: m_out<=8'b00001110;
        13'd416: m_out<=8'b00010101;
        13'd417: m_out<=8'b00011010;
        13'd418: m_out<=8'b11011101;
        13'd419: m_out<=8'b00000010;
        13'd420: m_out<=8'b11111001;
        13'd421: m_out<=8'b11110100;
        13'd422: m_out<=8'b11101100;
        13'd423: m_out<=8'b11011110;
        13'd424: m_out<=8'b00001100;
        13'd425: m_out<=8'b00011001;
        13'd426: m_out<=8'b00001011;
        13'd427: m_out<=8'b00010000;
        13'd428: m_out<=8'b11100100;
        13'd429: m_out<=8'b11100011;
        13'd430: m_out<=8'b00010010;
        13'd431: m_out<=8'b00000010;
        13'd432: m_out<=8'b01001001;
        13'd433: m_out<=8'b00000101;
        13'd434: m_out<=8'b00001000;
        13'd435: m_out<=8'b00001110;
        13'd436: m_out<=8'b11100101;
        13'd437: m_out<=8'b11110100;
        13'd438: m_out<=8'b00011000;
        13'd439: m_out<=8'b11110011;
        13'd440: m_out<=8'b11011111;
        13'd441: m_out<=8'b11101000;
        13'd442: m_out<=8'b11100110;
        13'd443: m_out<=8'b01000011;
        13'd444: m_out<=8'b11010110;
        13'd445: m_out<=8'b00000001;
        13'd446: m_out<=8'b00010111;
        13'd447: m_out<=8'b00010100;
        13'd448: m_out<=8'b00100100;
        13'd449: m_out<=8'b11111011;
        13'd450: m_out<=8'b00100111;
        13'd451: m_out<=8'b11111011;
        13'd452: m_out<=8'b00011011;
        13'd453: m_out<=8'b11101101;
        13'd454: m_out<=8'b00010000;
        13'd455: m_out<=8'b11110100;
        13'd456: m_out<=8'b11111111;
        13'd457: m_out<=8'b11001101;
        13'd458: m_out<=8'b00110011;
        13'd459: m_out<=8'b11010010;
        13'd460: m_out<=8'b00010110;
        13'd461: m_out<=8'b11101001;
        13'd462: m_out<=8'b11101100;
        13'd463: m_out<=8'b11111000;
        13'd464: m_out<=8'b00000010;
        13'd465: m_out<=8'b00001110;
        13'd466: m_out<=8'b11011101;
        13'd467: m_out<=8'b00010110;
        13'd468: m_out<=8'b11111000;
        13'd469: m_out<=8'b11101101;
        13'd470: m_out<=8'b00011110;
        13'd471: m_out<=8'b00011100;
        13'd472: m_out<=8'b11110011;
        13'd473: m_out<=8'b00001000;
        13'd474: m_out<=8'b00010100;
        13'd475: m_out<=8'b00010011;
        13'd476: m_out<=8'b00001000;
        13'd477: m_out<=8'b00001010;
        13'd478: m_out<=8'b00001111;
        13'd479: m_out<=8'b11110111;
        13'd480: m_out<=8'b00010010;
        13'd481: m_out<=8'b11111110;
        13'd482: m_out<=8'b00001100;
        13'd483: m_out<=8'b00011100;
        13'd484: m_out<=8'b11100100;
        13'd485: m_out<=8'b11100011;
        13'd486: m_out<=8'b11110100;
        13'd487: m_out<=8'b01000111;
        13'd488: m_out<=8'b11101110;
        13'd489: m_out<=8'b00001100;
        13'd490: m_out<=8'b00011011;
        13'd491: m_out<=8'b00101010;
        13'd492: m_out<=8'b00001010;
        13'd493: m_out<=8'b11111111;
        13'd494: m_out<=8'b11111011;
        13'd495: m_out<=8'b11000010;
        13'd496: m_out<=8'b00011111;
        13'd497: m_out<=8'b11011100;
        13'd498: m_out<=8'b00001000;
        13'd499: m_out<=8'b00010000;
        13'd500: m_out<=8'b00101001;
        13'd501: m_out<=8'b00011110;
        13'd502: m_out<=8'b11110010;
        13'd503: m_out<=8'b11111000;
        13'd504: m_out<=8'b10110010;
        13'd505: m_out<=8'b11110000;
        13'd506: m_out<=8'b00100010;
        13'd507: m_out<=8'b11100010;
        13'd508: m_out<=8'b00000010;
        13'd509: m_out<=8'b11100010;
        13'd510: m_out<=8'b11100110;
        13'd511: m_out<=8'b11011101;
        13'd512: m_out<=8'b00000001;
        13'd513: m_out<=8'b00011111;
        13'd514: m_out<=8'b00011000;
        13'd515: m_out<=8'b11111001;
        13'd516: m_out<=8'b00001100;
        13'd517: m_out<=8'b00010001;
        13'd518: m_out<=8'b11111000;
        13'd519: m_out<=8'b00000111;
        13'd520: m_out<=8'b11101111;
        13'd521: m_out<=8'b11111011;
        13'd522: m_out<=8'b11110111;
        13'd523: m_out<=8'b11101001;
        13'd524: m_out<=8'b11101100;
        13'd525: m_out<=8'b00011010;
        13'd526: m_out<=8'b00001100;
        13'd527: m_out<=8'b11101010;
        13'd528: m_out<=8'b11110011;
        13'd529: m_out<=8'b00011100;
        13'd530: m_out<=8'b11110011;
        13'd531: m_out<=8'b00111000;
        13'd532: m_out<=8'b11011101;
        13'd533: m_out<=8'b00000010;
        13'd534: m_out<=8'b00000101;
        13'd535: m_out<=8'b11100101;
        13'd536: m_out<=8'b11110001;
        13'd537: m_out<=8'b11011110;
        13'd538: m_out<=8'b11110011;
        13'd539: m_out<=8'b01001010;
        13'd540: m_out<=8'b00010101;
        13'd541: m_out<=8'b11111010;
        13'd542: m_out<=8'b00010010;
        13'd543: m_out<=8'b00010100;
        13'd544: m_out<=8'b11111000;
        13'd545: m_out<=8'b00001010;
        13'd546: m_out<=8'b11100111;
        13'd547: m_out<=8'b11110001;
        13'd548: m_out<=8'b11100100;
        13'd549: m_out<=8'b11100100;
        13'd550: m_out<=8'b11011100;
        13'd551: m_out<=8'b11110101;
        13'd552: m_out<=8'b11011111;
        13'd553: m_out<=8'b00000101;
        13'd554: m_out<=8'b11001101;
        13'd555: m_out<=8'b00100000;
        13'd556: m_out<=8'b00001011;
        13'd557: m_out<=8'b11011100;
        13'd558: m_out<=8'b00010110;
        13'd559: m_out<=8'b00001011;
        13'd560: m_out<=8'b00010001;
        13'd561: m_out<=8'b11101110;
        13'd562: m_out<=8'b11110111;
        13'd563: m_out<=8'b00000001;
        13'd564: m_out<=8'b11100001;
        13'd565: m_out<=8'b00000000;
        13'd566: m_out<=8'b00110001;
        13'd567: m_out<=8'b00001011;
        13'd568: m_out<=8'b11001111;
        13'd569: m_out<=8'b11101111;
        13'd570: m_out<=8'b00000001;
        13'd571: m_out<=8'b11100001;
        13'd572: m_out<=8'b11101001;
        13'd573: m_out<=8'b11100110;
        13'd574: m_out<=8'b11001011;
        13'd575: m_out<=8'b00001101;
        13'd576: m_out<=8'b00011110;
        13'd577: m_out<=8'b11110110;
        13'd578: m_out<=8'b00000010;
        13'd579: m_out<=8'b11110101;
        13'd580: m_out<=8'b00100001;
        13'd581: m_out<=8'b11011000;
        13'd582: m_out<=8'b11101001;
        13'd583: m_out<=8'b11111111;
        13'd584: m_out<=8'b00111101;
        13'd585: m_out<=8'b11111001;
        13'd586: m_out<=8'b00010000;
        13'd587: m_out<=8'b00100111;
        13'd588: m_out<=8'b00000000;
        13'd589: m_out<=8'b11100001;
        13'd590: m_out<=8'b00010000;
        13'd591: m_out<=8'b11010111;
        13'd592: m_out<=8'b11110100;
        13'd593: m_out<=8'b11101111;
        13'd594: m_out<=8'b00000110;
        13'd595: m_out<=8'b00100110;
        13'd596: m_out<=8'b00001110;
        13'd597: m_out<=8'b11100001;
        13'd598: m_out<=8'b00000111;
        13'd599: m_out<=8'b00010111;
        13'd600: m_out<=8'b00000001;
        13'd601: m_out<=8'b00010000;
        13'd602: m_out<=8'b00000101;
        13'd603: m_out<=8'b00000001;
        13'd604: m_out<=8'b00011101;
        13'd605: m_out<=8'b00010011;
        13'd606: m_out<=8'b11001110;
        13'd607: m_out<=8'b11101001;
        13'd608: m_out<=8'b00001110;
        13'd609: m_out<=8'b10111011;
        13'd610: m_out<=8'b11111011;
        13'd611: m_out<=8'b00000001;
        13'd612: m_out<=8'b00001010;
        13'd613: m_out<=8'b00000010;
        13'd614: m_out<=8'b00001011;
        13'd615: m_out<=8'b00010010;
        13'd616: m_out<=8'b11111100;
        13'd617: m_out<=8'b00011100;
        13'd618: m_out<=8'b00000111;
        13'd619: m_out<=8'b11110110;
        13'd620: m_out<=8'b11011100;
        13'd621: m_out<=8'b00011000;
        13'd622: m_out<=8'b00011001;
        13'd623: m_out<=8'b00110110;
        13'd624: m_out<=8'b00100111;
        13'd625: m_out<=8'b11101111;
        13'd626: m_out<=8'b00001011;
        13'd627: m_out<=8'b11011000;
        13'd628: m_out<=8'b11111011;
        13'd629: m_out<=8'b11101100;
        13'd630: m_out<=8'b11011010;
        13'd631: m_out<=8'b11111110;
        13'd632: m_out<=8'b11011101;
        13'd633: m_out<=8'b00011010;
        13'd634: m_out<=8'b11011110;
        13'd635: m_out<=8'b00010011;
        13'd636: m_out<=8'b00000010;
        13'd637: m_out<=8'b11100100;
        13'd638: m_out<=8'b00010101;
        13'd639: m_out<=8'b11111100;
        13'd640: m_out<=8'b00000101;
        13'd641: m_out<=8'b11110000;
        13'd642: m_out<=8'b00001111;
        13'd643: m_out<=8'b11110000;
        13'd644: m_out<=8'b00001100;
        13'd645: m_out<=8'b11101110;
        13'd646: m_out<=8'b00110011;
        13'd647: m_out<=8'b00011110;
        13'd648: m_out<=8'b11110011;
        13'd649: m_out<=8'b11111010;
        13'd650: m_out<=8'b11111100;
        13'd651: m_out<=8'b11101100;
        13'd652: m_out<=8'b11011110;
        13'd653: m_out<=8'b00010001;
        13'd654: m_out<=8'b00000101;
        13'd655: m_out<=8'b11110101;
        13'd656: m_out<=8'b11111001;
        13'd657: m_out<=8'b11101011;
        13'd658: m_out<=8'b00010101;
        13'd659: m_out<=8'b00010111;
        13'd660: m_out<=8'b11110000;
        13'd661: m_out<=8'b11100000;
        13'd662: m_out<=8'b00010011;
        13'd663: m_out<=8'b11011010;
        13'd664: m_out<=8'b00000011;
        13'd665: m_out<=8'b00011001;
        13'd666: m_out<=8'b00001110;
        13'd667: m_out<=8'b11011010;
        13'd668: m_out<=8'b11110110;
        13'd669: m_out<=8'b11110000;
        13'd670: m_out<=8'b11101100;
        13'd671: m_out<=8'b00011111;
        13'd672: m_out<=8'b11110001;
        13'd673: m_out<=8'b00100010;
        13'd674: m_out<=8'b00010000;
        13'd675: m_out<=8'b00110101;
        13'd676: m_out<=8'b00001000;
        13'd677: m_out<=8'b00001001;
        13'd678: m_out<=8'b11101010;
        13'd679: m_out<=8'b11100101;
        13'd680: m_out<=8'b11101101;
        13'd681: m_out<=8'b00101111;
        13'd682: m_out<=8'b00001001;
        13'd683: m_out<=8'b00000110;
        13'd684: m_out<=8'b11110101;
        13'd685: m_out<=8'b00100010;
        13'd686: m_out<=8'b11011011;
        13'd687: m_out<=8'b00000100;
        13'd688: m_out<=8'b11001010;
        13'd689: m_out<=8'b11111001;
        13'd690: m_out<=8'b11011100;
        13'd691: m_out<=8'b00010111;
        13'd692: m_out<=8'b11110010;
        13'd693: m_out<=8'b00000000;
        13'd694: m_out<=8'b11111101;
        13'd695: m_out<=8'b11011100;
        13'd696: m_out<=8'b11010010;
        13'd697: m_out<=8'b00001011;
        13'd698: m_out<=8'b00000101;
        13'd699: m_out<=8'b11101001;
        13'd700: m_out<=8'b11110000;
        13'd701: m_out<=8'b11110101;
        13'd702: m_out<=8'b00010100;
        13'd703: m_out<=8'b00101110;
        13'd704: m_out<=8'b00101011;
        13'd705: m_out<=8'b11110001;
        13'd706: m_out<=8'b00110000;
        13'd707: m_out<=8'b11110111;
        13'd708: m_out<=8'b11100011;
        13'd709: m_out<=8'b00000001;
        13'd710: m_out<=8'b11110001;
        13'd711: m_out<=8'b11011001;
        13'd712: m_out<=8'b11110001;
        13'd713: m_out<=8'b00001010;
        13'd714: m_out<=8'b00000100;
        13'd715: m_out<=8'b11110010;
        13'd716: m_out<=8'b00111101;
        13'd717: m_out<=8'b00110100;
        13'd718: m_out<=8'b00010000;
        13'd719: m_out<=8'b11011000;
        13'd720: m_out<=8'b00000110;
        13'd721: m_out<=8'b00000011;
        13'd722: m_out<=8'b00000000;
        13'd723: m_out<=8'b00000110;
        13'd724: m_out<=8'b11110010;
        13'd725: m_out<=8'b11111001;
        13'd726: m_out<=8'b11101000;
        13'd727: m_out<=8'b11101000;
        13'd728: m_out<=8'b11010101;
        13'd729: m_out<=8'b00011100;
        13'd730: m_out<=8'b11010110;
        13'd731: m_out<=8'b00010100;
        13'd732: m_out<=8'b00011010;
        13'd733: m_out<=8'b00001011;
        13'd734: m_out<=8'b00000010;
        13'd735: m_out<=8'b11100101;
        13'd736: m_out<=8'b10111101;
        13'd737: m_out<=8'b00000100;
        13'd738: m_out<=8'b00001101;
        13'd739: m_out<=8'b11100010;
        13'd740: m_out<=8'b11000110;
        13'd741: m_out<=8'b11110101;
        13'd742: m_out<=8'b11110010;
        13'd743: m_out<=8'b11110100;
        13'd744: m_out<=8'b00011110;
        13'd745: m_out<=8'b11110011;
        13'd746: m_out<=8'b00011010;
        13'd747: m_out<=8'b00000101;
        13'd748: m_out<=8'b11101101;
        13'd749: m_out<=8'b11100100;
        13'd750: m_out<=8'b11101100;
        13'd751: m_out<=8'b00011100;
        13'd752: m_out<=8'b11100111;
        13'd753: m_out<=8'b11100111;
        13'd754: m_out<=8'b11011111;
        13'd755: m_out<=8'b11111101;
        13'd756: m_out<=8'b11110110;
        13'd757: m_out<=8'b11100101;
        13'd758: m_out<=8'b00010110;
        13'd759: m_out<=8'b11101011;
        13'd760: m_out<=8'b11111011;
        13'd761: m_out<=8'b00011110;
        13'd762: m_out<=8'b00011010;
        13'd763: m_out<=8'b00000100;
        13'd764: m_out<=8'b11101101;
        13'd765: m_out<=8'b11110010;
        13'd766: m_out<=8'b11110001;
        13'd767: m_out<=8'b11111010;
        13'd768: m_out<=8'b00011000;
        13'd769: m_out<=8'b00001100;
        13'd770: m_out<=8'b00000011;
        13'd771: m_out<=8'b11110011;
        13'd772: m_out<=8'b11111111;
        13'd773: m_out<=8'b00010011;
        13'd774: m_out<=8'b00000011;
        13'd775: m_out<=8'b11110011;
        13'd776: m_out<=8'b00001101;
        13'd777: m_out<=8'b11011000;
        13'd778: m_out<=8'b11101000;
        13'd779: m_out<=8'b00000000;
        13'd780: m_out<=8'b11101110;
        13'd781: m_out<=8'b11001110;
        13'd782: m_out<=8'b11110000;
        13'd783: m_out<=8'b00011101;
        13'd784: m_out<=8'b00010011;
        13'd785: m_out<=8'b00001110;
        13'd786: m_out<=8'b00010001;
        13'd787: m_out<=8'b11111001;
        13'd788: m_out<=8'b00010100;
        13'd789: m_out<=8'b00001111;
        13'd790: m_out<=8'b11101011;
        13'd791: m_out<=8'b11111110;
        13'd792: m_out<=8'b00000101;
        13'd793: m_out<=8'b00101100;
        13'd794: m_out<=8'b11110101;
        13'd795: m_out<=8'b11111011;
        13'd796: m_out<=8'b11101000;
        13'd797: m_out<=8'b00101110;
        13'd798: m_out<=8'b00100001;
        13'd799: m_out<=8'b11110011;
        13'd800: m_out<=8'b00001101;
        13'd801: m_out<=8'b00100111;
        13'd802: m_out<=8'b00001101;
        13'd803: m_out<=8'b11111000;
        13'd804: m_out<=8'b00101100;
        13'd805: m_out<=8'b11011110;
        13'd806: m_out<=8'b00100110;
        13'd807: m_out<=8'b11110110;
        13'd808: m_out<=8'b00001100;
        13'd809: m_out<=8'b00001110;
        13'd810: m_out<=8'b00110000;
        13'd811: m_out<=8'b11010100;
        13'd812: m_out<=8'b00001000;
        13'd813: m_out<=8'b11101111;
        13'd814: m_out<=8'b11110100;
        13'd815: m_out<=8'b11110001;
        13'd816: m_out<=8'b11010011;
        13'd817: m_out<=8'b11110001;
        13'd818: m_out<=8'b11100001;
        13'd819: m_out<=8'b11100100;
        13'd820: m_out<=8'b11111000;
        13'd821: m_out<=8'b11110011;
        13'd822: m_out<=8'b00000100;
        13'd823: m_out<=8'b00000001;
        13'd824: m_out<=8'b00100011;
        13'd825: m_out<=8'b00000100;
        13'd826: m_out<=8'b11011100;
        13'd827: m_out<=8'b00001101;
        13'd828: m_out<=8'b11111010;
        13'd829: m_out<=8'b11010101;
        13'd830: m_out<=8'b00000001;
        13'd831: m_out<=8'b00001010;
        13'd832: m_out<=8'b11110111;
        13'd833: m_out<=8'b11100011;
        13'd834: m_out<=8'b00010000;
        13'd835: m_out<=8'b00001101;
        13'd836: m_out<=8'b00000100;
        13'd837: m_out<=8'b00000100;
        13'd838: m_out<=8'b00011011;
        13'd839: m_out<=8'b00000111;
        13'd840: m_out<=8'b11101101;
        13'd841: m_out<=8'b01001100;
        13'd842: m_out<=8'b00001011;
        13'd843: m_out<=8'b00000101;
        13'd844: m_out<=8'b00001100;
        13'd845: m_out<=8'b00011010;
        13'd846: m_out<=8'b00001000;
        13'd847: m_out<=8'b00011010;
        13'd848: m_out<=8'b00111111;
        13'd849: m_out<=8'b11101001;
        13'd850: m_out<=8'b00100001;
        13'd851: m_out<=8'b00001000;
        13'd852: m_out<=8'b11111001;
        13'd853: m_out<=8'b00010111;
        13'd854: m_out<=8'b11110100;
        13'd855: m_out<=8'b00011010;
        13'd856: m_out<=8'b11111111;
        13'd857: m_out<=8'b00000110;
        13'd858: m_out<=8'b10110110;
        13'd859: m_out<=8'b00000000;
        13'd860: m_out<=8'b11111101;
        13'd861: m_out<=8'b11101101;
        13'd862: m_out<=8'b11011010;
        13'd863: m_out<=8'b11111101;
        13'd864: m_out<=8'b00101100;
        13'd865: m_out<=8'b00001011;
        13'd866: m_out<=8'b11111110;
        13'd867: m_out<=8'b11100111;
        13'd868: m_out<=8'b00100111;
        13'd869: m_out<=8'b00010101;
        13'd870: m_out<=8'b00011011;
        13'd871: m_out<=8'b11110011;
        13'd872: m_out<=8'b00100001;
        13'd873: m_out<=8'b00011010;
        13'd874: m_out<=8'b11110110;
        13'd875: m_out<=8'b00000010;
        13'd876: m_out<=8'b11111010;
        13'd877: m_out<=8'b11111110;
        13'd878: m_out<=8'b00011111;
        13'd879: m_out<=8'b11111001;
        13'd880: m_out<=8'b11111111;
        13'd881: m_out<=8'b11111111;
        13'd882: m_out<=8'b00000001;
        13'd883: m_out<=8'b11101011;
        13'd884: m_out<=8'b00000010;
        13'd885: m_out<=8'b00000010;
        13'd886: m_out<=8'b11100011;
        13'd887: m_out<=8'b00010000;
        13'd888: m_out<=8'b00001011;
        13'd889: m_out<=8'b00100100;
        13'd890: m_out<=8'b11100101;
        13'd891: m_out<=8'b11111110;
        13'd892: m_out<=8'b11010101;
        13'd893: m_out<=8'b00010000;
        13'd894: m_out<=8'b11000111;
        13'd895: m_out<=8'b00001101;
        13'd896: m_out<=8'b00011010;
        13'd897: m_out<=8'b11110000;
        13'd898: m_out<=8'b00011101;
        13'd899: m_out<=8'b11101101;
        13'd900: m_out<=8'b00011111;
        13'd901: m_out<=8'b00000000;
        13'd902: m_out<=8'b00101100;
        13'd903: m_out<=8'b11011010;
        13'd904: m_out<=8'b00011111;
        13'd905: m_out<=8'b11101100;
        13'd906: m_out<=8'b11111111;
        13'd907: m_out<=8'b00001000;
        13'd908: m_out<=8'b11110111;
        13'd909: m_out<=8'b00011000;
        13'd910: m_out<=8'b00010111;
        13'd911: m_out<=8'b00000010;
        13'd912: m_out<=8'b11111110;
        13'd913: m_out<=8'b00100000;
        13'd914: m_out<=8'b00101010;
        13'd915: m_out<=8'b11111100;
        13'd916: m_out<=8'b11010111;
        13'd917: m_out<=8'b00000010;
        13'd918: m_out<=8'b11111101;
        13'd919: m_out<=8'b00100101;
        13'd920: m_out<=8'b11110111;
        13'd921: m_out<=8'b11101110;
        13'd922: m_out<=8'b11101100;
        13'd923: m_out<=8'b11101011;
        13'd924: m_out<=8'b00010010;
        13'd925: m_out<=8'b11010111;
        13'd926: m_out<=8'b11101011;
        13'd927: m_out<=8'b11110100;
        13'd928: m_out<=8'b00000101;
        13'd929: m_out<=8'b00011111;
        13'd930: m_out<=8'b01001011;
        13'd931: m_out<=8'b11111111;
        13'd932: m_out<=8'b11100111;
        13'd933: m_out<=8'b11111001;
        13'd934: m_out<=8'b11110011;
        13'd935: m_out<=8'b11110111;
        13'd936: m_out<=8'b00000000;
        13'd937: m_out<=8'b00001010;
        13'd938: m_out<=8'b11011100;
        13'd939: m_out<=8'b11101101;
        13'd940: m_out<=8'b11101000;
        13'd941: m_out<=8'b00011010;
        13'd942: m_out<=8'b00010111;
        13'd943: m_out<=8'b00001010;
        13'd944: m_out<=8'b11100100;
        13'd945: m_out<=8'b00000011;
        13'd946: m_out<=8'b11111011;
        13'd947: m_out<=8'b00001111;
        13'd948: m_out<=8'b11011101;
        13'd949: m_out<=8'b11101011;
        13'd950: m_out<=8'b00010011;
        13'd951: m_out<=8'b11110101;
        13'd952: m_out<=8'b11110010;
        13'd953: m_out<=8'b00000010;
        13'd954: m_out<=8'b00000101;
        13'd955: m_out<=8'b00101110;
        13'd956: m_out<=8'b11011011;
        13'd957: m_out<=8'b11101011;
        13'd958: m_out<=8'b11010001;
        13'd959: m_out<=8'b00011110;
        13'd960: m_out<=8'b11011101;
        13'd961: m_out<=8'b00110011;
        13'd962: m_out<=8'b11101110;
        13'd963: m_out<=8'b00101101;
        13'd964: m_out<=8'b11101011;
        13'd965: m_out<=8'b11011111;
        13'd966: m_out<=8'b11111000;
        13'd967: m_out<=8'b11011110;
        13'd968: m_out<=8'b11111011;
        13'd969: m_out<=8'b00000001;
        13'd970: m_out<=8'b00000110;
        13'd971: m_out<=8'b11111101;
        13'd972: m_out<=8'b11110000;
        13'd973: m_out<=8'b11111101;
        13'd974: m_out<=8'b00001000;
        13'd975: m_out<=8'b00010000;
        13'd976: m_out<=8'b11101111;
        13'd977: m_out<=8'b11110111;
        13'd978: m_out<=8'b11111000;
        13'd979: m_out<=8'b11010100;
        13'd980: m_out<=8'b11100011;
        13'd981: m_out<=8'b00000111;
        13'd982: m_out<=8'b00100001;
        13'd983: m_out<=8'b00000010;
        13'd984: m_out<=8'b00100001;
        13'd985: m_out<=8'b11100000;
        13'd986: m_out<=8'b00000011;
        13'd987: m_out<=8'b00001011;
        13'd988: m_out<=8'b00010000;
        13'd989: m_out<=8'b00011010;
        13'd990: m_out<=8'b00010001;
        13'd991: m_out<=8'b00001011;
        13'd992: m_out<=8'b00010010;
        13'd993: m_out<=8'b11101101;
        13'd994: m_out<=8'b11100000;
        13'd995: m_out<=8'b11110010;
        13'd996: m_out<=8'b00010111;
        13'd997: m_out<=8'b00001111;
        13'd998: m_out<=8'b11010110;
        13'd999: m_out<=8'b00000000;
        13'd1000: m_out<=8'b11101100;
        13'd1001: m_out<=8'b11101111;
        13'd1002: m_out<=8'b00001010;
        13'd1003: m_out<=8'b11101110;
        13'd1004: m_out<=8'b11101000;
        13'd1005: m_out<=8'b00000111;
        13'd1006: m_out<=8'b00100100;
        13'd1007: m_out<=8'b11100001;
        13'd1008: m_out<=8'b00000101;
        13'd1009: m_out<=8'b00001111;
        13'd1010: m_out<=8'b00011001;
        13'd1011: m_out<=8'b11101010;
        13'd1012: m_out<=8'b11100011;
        13'd1013: m_out<=8'b00010001;
        13'd1014: m_out<=8'b01001001;
        13'd1015: m_out<=8'b00000001;
        13'd1016: m_out<=8'b11111101;
        13'd1017: m_out<=8'b11111011;
        13'd1018: m_out<=8'b00101011;
        13'd1019: m_out<=8'b11010001;
        13'd1020: m_out<=8'b00100000;
        13'd1021: m_out<=8'b11110001;
        13'd1022: m_out<=8'b00100001;
        13'd1023: m_out<=8'b00000010;
        13'd1024: m_out<=8'b11010101;
        13'd1025: m_out<=8'b00001011;
        13'd1026: m_out<=8'b00000111;
        13'd1027: m_out<=8'b00001111;
        13'd1028: m_out<=8'b11110110;
        13'd1029: m_out<=8'b11101111;
        13'd1030: m_out<=8'b00001011;
        13'd1031: m_out<=8'b00011000;
        13'd1032: m_out<=8'b11111111;
        13'd1033: m_out<=8'b11111010;
        13'd1034: m_out<=8'b11100011;
        13'd1035: m_out<=8'b11100111;
        13'd1036: m_out<=8'b00001010;
        13'd1037: m_out<=8'b00000011;
        13'd1038: m_out<=8'b00011110;
        13'd1039: m_out<=8'b11101010;
        13'd1040: m_out<=8'b11101001;
        13'd1041: m_out<=8'b00010010;
        13'd1042: m_out<=8'b11101101;
        13'd1043: m_out<=8'b11110001;
        13'd1044: m_out<=8'b00100100;
        13'd1045: m_out<=8'b11101100;
        13'd1046: m_out<=8'b00000101;
        13'd1047: m_out<=8'b11111000;
        13'd1048: m_out<=8'b00111100;
        13'd1049: m_out<=8'b11110010;
        13'd1050: m_out<=8'b00000001;
        13'd1051: m_out<=8'b11110111;
        13'd1052: m_out<=8'b00001001;
        13'd1053: m_out<=8'b11101010;
        13'd1054: m_out<=8'b00011001;
        13'd1055: m_out<=8'b11111110;
        13'd1056: m_out<=8'b00010010;
        13'd1057: m_out<=8'b11100111;
        13'd1058: m_out<=8'b00010011;
        13'd1059: m_out<=8'b11100110;
        13'd1060: m_out<=8'b00010100;
        13'd1061: m_out<=8'b00000111;
        13'd1062: m_out<=8'b11100010;
        13'd1063: m_out<=8'b11101101;
        13'd1064: m_out<=8'b00100111;
        13'd1065: m_out<=8'b11111100;
        13'd1066: m_out<=8'b00001001;
        13'd1067: m_out<=8'b00011100;
        13'd1068: m_out<=8'b00010001;
        13'd1069: m_out<=8'b11101010;
        13'd1070: m_out<=8'b00001101;
        13'd1071: m_out<=8'b11100000;
        13'd1072: m_out<=8'b11011101;
        13'd1073: m_out<=8'b11101110;
        13'd1074: m_out<=8'b11100110;
        13'd1075: m_out<=8'b00000101;
        13'd1076: m_out<=8'b11101110;
        13'd1077: m_out<=8'b00000110;
        13'd1078: m_out<=8'b11110011;
        13'd1079: m_out<=8'b11101110;
        13'd1080: m_out<=8'b11010010;
        13'd1081: m_out<=8'b00000000;
        13'd1082: m_out<=8'b00100010;
        13'd1083: m_out<=8'b11110110;
        13'd1084: m_out<=8'b00000010;
        13'd1085: m_out<=8'b11111110;
        13'd1086: m_out<=8'b00100000;
        13'd1087: m_out<=8'b11101110;
        13'd1088: m_out<=8'b00000100;
        13'd1089: m_out<=8'b11101011;
        13'd1090: m_out<=8'b00010010;
        13'd1091: m_out<=8'b11001100;
        13'd1092: m_out<=8'b00000100;
        13'd1093: m_out<=8'b00110110;
        13'd1094: m_out<=8'b11111110;
        13'd1095: m_out<=8'b00110101;
        13'd1096: m_out<=8'b11111001;
        13'd1097: m_out<=8'b11111000;
        13'd1098: m_out<=8'b00010100;
        13'd1099: m_out<=8'b00100101;
        13'd1100: m_out<=8'b11110010;
        13'd1101: m_out<=8'b11011111;
        13'd1102: m_out<=8'b00011110;
        13'd1103: m_out<=8'b00101000;
        13'd1104: m_out<=8'b00001101;
        13'd1105: m_out<=8'b00011000;
        13'd1106: m_out<=8'b11100011;
        13'd1107: m_out<=8'b00010110;
        13'd1108: m_out<=8'b11111010;
        13'd1109: m_out<=8'b11001100;
        13'd1110: m_out<=8'b11100111;
        13'd1111: m_out<=8'b00010001;
        13'd1112: m_out<=8'b11011001;
        13'd1113: m_out<=8'b11111110;
        13'd1114: m_out<=8'b11111000;
        13'd1115: m_out<=8'b11110100;
        13'd1116: m_out<=8'b00010101;
        13'd1117: m_out<=8'b11111011;
        13'd1118: m_out<=8'b11111111;
        13'd1119: m_out<=8'b00101001;
        13'd1120: m_out<=8'b11111100;
        13'd1121: m_out<=8'b00010110;
        13'd1122: m_out<=8'b11100000;
        13'd1123: m_out<=8'b00001011;
        13'd1124: m_out<=8'b11100010;
        13'd1125: m_out<=8'b11100010;
        13'd1126: m_out<=8'b11111000;
        13'd1127: m_out<=8'b00001010;
        13'd1128: m_out<=8'b11101000;
        13'd1129: m_out<=8'b00000111;
        13'd1130: m_out<=8'b11110000;
        13'd1131: m_out<=8'b00010000;
        13'd1132: m_out<=8'b00001000;
        13'd1133: m_out<=8'b11111100;
        13'd1134: m_out<=8'b11111001;
        13'd1135: m_out<=8'b11111000;
        13'd1136: m_out<=8'b00100001;
        13'd1137: m_out<=8'b11101111;
        13'd1138: m_out<=8'b11101000;
        13'd1139: m_out<=8'b11101011;
        13'd1140: m_out<=8'b11011011;
        13'd1141: m_out<=8'b00010011;
        13'd1142: m_out<=8'b00001111;
        13'd1143: m_out<=8'b00011110;
        13'd1144: m_out<=8'b11101001;
        13'd1145: m_out<=8'b11111101;
        13'd1146: m_out<=8'b11111000;
        13'd1147: m_out<=8'b11110100;
        13'd1148: m_out<=8'b11101010;
        13'd1149: m_out<=8'b00001011;
        13'd1150: m_out<=8'b11110111;
        13'd1151: m_out<=8'b11110011;
        13'd1152: m_out<=8'b11011010;
        13'd1153: m_out<=8'b11110110;
        13'd1154: m_out<=8'b00011001;
        13'd1155: m_out<=8'b00100000;
        13'd1156: m_out<=8'b11111111;
        13'd1157: m_out<=8'b00100100;
        13'd1158: m_out<=8'b11111000;
        13'd1159: m_out<=8'b00000100;
        13'd1160: m_out<=8'b00011000;
        13'd1161: m_out<=8'b11101001;
        13'd1162: m_out<=8'b00001001;
        13'd1163: m_out<=8'b00101100;
        13'd1164: m_out<=8'b11000101;
        13'd1165: m_out<=8'b00010011;
        13'd1166: m_out<=8'b00011010;
        13'd1167: m_out<=8'b00001111;
        13'd1168: m_out<=8'b00100100;
        13'd1169: m_out<=8'b00011000;
        13'd1170: m_out<=8'b11101010;
        13'd1171: m_out<=8'b00101111;
        13'd1172: m_out<=8'b00010110;
        13'd1173: m_out<=8'b11011011;
        13'd1174: m_out<=8'b11111110;
        13'd1175: m_out<=8'b00100000;
        13'd1176: m_out<=8'b11111010;
        13'd1177: m_out<=8'b00000100;
        13'd1178: m_out<=8'b11101110;
        13'd1179: m_out<=8'b11110111;
        13'd1180: m_out<=8'b00000111;
        13'd1181: m_out<=8'b11100111;
        13'd1182: m_out<=8'b11001100;
        13'd1183: m_out<=8'b00011001;
        13'd1184: m_out<=8'b11101010;
        13'd1185: m_out<=8'b00000001;
        13'd1186: m_out<=8'b11110111;
        13'd1187: m_out<=8'b11110000;
        13'd1188: m_out<=8'b11111011;
        13'd1189: m_out<=8'b11110000;
        13'd1190: m_out<=8'b00001000;
        13'd1191: m_out<=8'b11111010;
        13'd1192: m_out<=8'b11110101;
        13'd1193: m_out<=8'b11111110;
        13'd1194: m_out<=8'b00010001;
        13'd1195: m_out<=8'b11101001;
        13'd1196: m_out<=8'b11110100;
        13'd1197: m_out<=8'b00010101;
        13'd1198: m_out<=8'b00100010;
        13'd1199: m_out<=8'b11101001;
        13'd1200: m_out<=8'b00000011;
        13'd1201: m_out<=8'b11100010;
        13'd1202: m_out<=8'b11011011;
        13'd1203: m_out<=8'b11100100;
        13'd1204: m_out<=8'b11001111;
        13'd1205: m_out<=8'b11111000;
        13'd1206: m_out<=8'b11010001;
        13'd1207: m_out<=8'b11111100;
        13'd1208: m_out<=8'b11110010;
        13'd1209: m_out<=8'b00010010;
        13'd1210: m_out<=8'b00001110;
        13'd1211: m_out<=8'b11111011;
        13'd1212: m_out<=8'b00110011;
        13'd1213: m_out<=8'b11101000;
        13'd1214: m_out<=8'b00010010;
        13'd1215: m_out<=8'b11110001;
        13'd1216: m_out<=8'b00001011;
        13'd1217: m_out<=8'b11110100;
        13'd1218: m_out<=8'b11100110;
        13'd1219: m_out<=8'b11100010;
        13'd1220: m_out<=8'b00000010;
        13'd1221: m_out<=8'b00100100;
        13'd1222: m_out<=8'b11111001;
        13'd1223: m_out<=8'b11000110;
        13'd1224: m_out<=8'b11111010;
        13'd1225: m_out<=8'b00000001;
        13'd1226: m_out<=8'b11011101;
        13'd1227: m_out<=8'b00010010;
        13'd1228: m_out<=8'b00001110;
        13'd1229: m_out<=8'b00011111;
        13'd1230: m_out<=8'b00001010;
        13'd1231: m_out<=8'b00001010;
        13'd1232: m_out<=8'b00010100;
        13'd1233: m_out<=8'b00101101;
        13'd1234: m_out<=8'b11111101;
        13'd1235: m_out<=8'b00011111;
        13'd1236: m_out<=8'b00001111;
        13'd1237: m_out<=8'b11110101;
        13'd1238: m_out<=8'b00011000;
        13'd1239: m_out<=8'b00010000;
        13'd1240: m_out<=8'b11110001;
        13'd1241: m_out<=8'b11110101;
        13'd1242: m_out<=8'b00000000;
        13'd1243: m_out<=8'b11111100;
        13'd1244: m_out<=8'b00001110;
        13'd1245: m_out<=8'b00010111;
        13'd1246: m_out<=8'b11110100;
        13'd1247: m_out<=8'b11000111;
        13'd1248: m_out<=8'b11100001;
        13'd1249: m_out<=8'b01010101;
        13'd1250: m_out<=8'b11111101;
        13'd1251: m_out<=8'b11110000;
        13'd1252: m_out<=8'b00001011;
        13'd1253: m_out<=8'b00001110;
        13'd1254: m_out<=8'b00010100;
        13'd1255: m_out<=8'b00001001;
        13'd1256: m_out<=8'b11101000;
        13'd1257: m_out<=8'b11101100;
        13'd1258: m_out<=8'b00100000;
        13'd1259: m_out<=8'b00000101;
        13'd1260: m_out<=8'b00000000;
        13'd1261: m_out<=8'b00010100;
        13'd1262: m_out<=8'b00010101;
        13'd1263: m_out<=8'b11001111;
        13'd1264: m_out<=8'b00000100;
        13'd1265: m_out<=8'b11110000;
        13'd1266: m_out<=8'b00011101;
        13'd1267: m_out<=8'b11110001;
        13'd1268: m_out<=8'b11110000;
        13'd1269: m_out<=8'b11010011;
        13'd1270: m_out<=8'b11000100;
        13'd1271: m_out<=8'b00000100;
        13'd1272: m_out<=8'b11111100;
        13'd1273: m_out<=8'b00011000;
        13'd1274: m_out<=8'b00000111;
        13'd1275: m_out<=8'b00000111;
        13'd1276: m_out<=8'b11011100;
        13'd1277: m_out<=8'b11100110;
        13'd1278: m_out<=8'b00010110;
        13'd1279: m_out<=8'b11101110;
        13'd1280: m_out<=8'b11101111;
        13'd1281: m_out<=8'b11111011;
        13'd1282: m_out<=8'b11111100;
        13'd1283: m_out<=8'b01000001;
        13'd1284: m_out<=8'b00001111;
        13'd1285: m_out<=8'b11010010;
        13'd1286: m_out<=8'b11001101;
        13'd1287: m_out<=8'b11100010;
        13'd1288: m_out<=8'b00000001;
        13'd1289: m_out<=8'b00010000;
        13'd1290: m_out<=8'b00001010;
        13'd1291: m_out<=8'b11111110;
        13'd1292: m_out<=8'b11110110;
        13'd1293: m_out<=8'b00101000;
        13'd1294: m_out<=8'b00000010;
        13'd1295: m_out<=8'b11100111;
        13'd1296: m_out<=8'b10110001;
        13'd1297: m_out<=8'b00010011;
        13'd1298: m_out<=8'b11111111;
        13'd1299: m_out<=8'b00010101;
        13'd1300: m_out<=8'b00010001;
        13'd1301: m_out<=8'b11001111;
        13'd1302: m_out<=8'b11111000;
        13'd1303: m_out<=8'b00000001;
        13'd1304: m_out<=8'b00011001;
        13'd1305: m_out<=8'b00000011;
        13'd1306: m_out<=8'b11111110;
        13'd1307: m_out<=8'b11100000;
        13'd1308: m_out<=8'b11111111;
        13'd1309: m_out<=8'b11010011;
        13'd1310: m_out<=8'b11110000;
        13'd1311: m_out<=8'b11011011;
        13'd1312: m_out<=8'b00100001;
        13'd1313: m_out<=8'b11111111;
        13'd1314: m_out<=8'b11110001;
        13'd1315: m_out<=8'b00010000;
        13'd1316: m_out<=8'b00101101;
        13'd1317: m_out<=8'b00001011;
        13'd1318: m_out<=8'b00100001;
        13'd1319: m_out<=8'b11100110;
        13'd1320: m_out<=8'b11101100;
        13'd1321: m_out<=8'b00010011;
        13'd1322: m_out<=8'b00110001;
        13'd1323: m_out<=8'b11100101;
        13'd1324: m_out<=8'b11110000;
        13'd1325: m_out<=8'b11111000;
        13'd1326: m_out<=8'b00011000;
        13'd1327: m_out<=8'b11111001;
        13'd1328: m_out<=8'b01000010;
        13'd1329: m_out<=8'b11111110;
        13'd1330: m_out<=8'b00010101;
        13'd1331: m_out<=8'b00010101;
        13'd1332: m_out<=8'b11111100;
        13'd1333: m_out<=8'b11101111;
        13'd1334: m_out<=8'b00000100;
        13'd1335: m_out<=8'b00001010;
        13'd1336: m_out<=8'b11011100;
        13'd1337: m_out<=8'b11101001;
        13'd1338: m_out<=8'b00001011;
        13'd1339: m_out<=8'b11110011;
        13'd1340: m_out<=8'b11101000;
        13'd1341: m_out<=8'b11110101;
        13'd1342: m_out<=8'b00000001;
        13'd1343: m_out<=8'b00101110;
        13'd1344: m_out<=8'b11110110;
        13'd1345: m_out<=8'b00000011;
        13'd1346: m_out<=8'b00010011;
        13'd1347: m_out<=8'b00001001;
        13'd1348: m_out<=8'b00001100;
        13'd1349: m_out<=8'b11111000;
        13'd1350: m_out<=8'b10110001;
        13'd1351: m_out<=8'b11110111;
        13'd1352: m_out<=8'b00000010;
        13'd1353: m_out<=8'b00001010;
        13'd1354: m_out<=8'b00011010;
        13'd1355: m_out<=8'b00011110;
        13'd1356: m_out<=8'b11111111;
        13'd1357: m_out<=8'b00000001;
        13'd1358: m_out<=8'b00100100;
        13'd1359: m_out<=8'b11100111;
        13'd1360: m_out<=8'b00101011;
        13'd1361: m_out<=8'b00001110;
        13'd1362: m_out<=8'b11111110;
        13'd1363: m_out<=8'b11110010;
        13'd1364: m_out<=8'b11101111;
        13'd1365: m_out<=8'b11101001;
        13'd1366: m_out<=8'b00010011;
        13'd1367: m_out<=8'b11001011;
        13'd1368: m_out<=8'b11101111;
        13'd1369: m_out<=8'b00010100;
        13'd1370: m_out<=8'b11110000;
        13'd1371: m_out<=8'b11111001;
        13'd1372: m_out<=8'b00010000;
        13'd1373: m_out<=8'b00000000;
        13'd1374: m_out<=8'b11111011;
        13'd1375: m_out<=8'b00100000;
        13'd1376: m_out<=8'b11000001;
        13'd1377: m_out<=8'b00001011;
        13'd1378: m_out<=8'b11110001;
        13'd1379: m_out<=8'b11101011;
        13'd1380: m_out<=8'b11110010;
        13'd1381: m_out<=8'b11111001;
        13'd1382: m_out<=8'b11101100;
        13'd1383: m_out<=8'b11111100;
        13'd1384: m_out<=8'b00001001;
        13'd1385: m_out<=8'b11110111;
        13'd1386: m_out<=8'b11110100;
        13'd1387: m_out<=8'b11111000;
        13'd1388: m_out<=8'b00001100;
        13'd1389: m_out<=8'b00101001;
        13'd1390: m_out<=8'b11111101;
        13'd1391: m_out<=8'b00101100;
        13'd1392: m_out<=8'b00100110;
        13'd1393: m_out<=8'b11111011;
        13'd1394: m_out<=8'b11111001;
        13'd1395: m_out<=8'b11101001;
        13'd1396: m_out<=8'b00010111;
        13'd1397: m_out<=8'b00011011;
        13'd1398: m_out<=8'b11011000;
        13'd1399: m_out<=8'b00010111;
        13'd1400: m_out<=8'b11111001;
        13'd1401: m_out<=8'b11100101;
        13'd1402: m_out<=8'b00001110;
        13'd1403: m_out<=8'b11110110;
        13'd1404: m_out<=8'b11111000;
        13'd1405: m_out<=8'b11101011;
        13'd1406: m_out<=8'b00100010;
        13'd1407: m_out<=8'b00100011;
        13'd1408: m_out<=8'b11111011;
        13'd1409: m_out<=8'b00001101;
        13'd1410: m_out<=8'b00001100;
        13'd1411: m_out<=8'b11100101;
        13'd1412: m_out<=8'b11110111;
        13'd1413: m_out<=8'b00000100;
        13'd1414: m_out<=8'b11101010;
        13'd1415: m_out<=8'b00110000;
        13'd1416: m_out<=8'b11111001;
        13'd1417: m_out<=8'b11100011;
        13'd1418: m_out<=8'b00010110;
        13'd1419: m_out<=8'b11111100;
        13'd1420: m_out<=8'b11100100;
        13'd1421: m_out<=8'b00011101;
        13'd1422: m_out<=8'b11100101;
        13'd1423: m_out<=8'b00011001;
        13'd1424: m_out<=8'b11111100;
        13'd1425: m_out<=8'b11110011;
        13'd1426: m_out<=8'b00000010;
        13'd1427: m_out<=8'b00000010;
        13'd1428: m_out<=8'b00000111;
        13'd1429: m_out<=8'b11101110;
        13'd1430: m_out<=8'b11100110;
        13'd1431: m_out<=8'b00000010;
        13'd1432: m_out<=8'b00100010;
        13'd1433: m_out<=8'b11100101;
        13'd1434: m_out<=8'b11101110;
        13'd1435: m_out<=8'b00001101;
        13'd1436: m_out<=8'b11010001;
        13'd1437: m_out<=8'b00000000;
        13'd1438: m_out<=8'b11011001;
        13'd1439: m_out<=8'b11100111;
        13'd1440: m_out<=8'b00001100;
        13'd1441: m_out<=8'b00000100;
        13'd1442: m_out<=8'b00101001;
        13'd1443: m_out<=8'b00000110;
        13'd1444: m_out<=8'b11110011;
        13'd1445: m_out<=8'b11101110;
        13'd1446: m_out<=8'b11110001;
        13'd1447: m_out<=8'b00011100;
        13'd1448: m_out<=8'b00101110;
        13'd1449: m_out<=8'b00011010;
        13'd1450: m_out<=8'b11111100;
        13'd1451: m_out<=8'b00010000;
        13'd1452: m_out<=8'b00001001;
        13'd1453: m_out<=8'b00100100;
        13'd1454: m_out<=8'b11111011;
        13'd1455: m_out<=8'b11101111;
        13'd1456: m_out<=8'b00100100;
        13'd1457: m_out<=8'b11100111;
        13'd1458: m_out<=8'b00110011;
        13'd1459: m_out<=8'b11011011;
        13'd1460: m_out<=8'b00101001;
        13'd1461: m_out<=8'b00000010;
        13'd1462: m_out<=8'b00011100;
        13'd1463: m_out<=8'b11110101;
        13'd1464: m_out<=8'b11010110;
        13'd1465: m_out<=8'b11011000;
        13'd1466: m_out<=8'b00011001;
        13'd1467: m_out<=8'b00010100;
        13'd1468: m_out<=8'b11001100;
        13'd1469: m_out<=8'b11111000;
        13'd1470: m_out<=8'b00001001;
        13'd1471: m_out<=8'b00101011;
        13'd1472: m_out<=8'b00011100;
        13'd1473: m_out<=8'b11100100;
        13'd1474: m_out<=8'b00001011;
        13'd1475: m_out<=8'b00000101;
        13'd1476: m_out<=8'b00000010;
        13'd1477: m_out<=8'b11101011;
        13'd1478: m_out<=8'b00000110;
        13'd1479: m_out<=8'b11111010;
        13'd1480: m_out<=8'b00011001;
        13'd1481: m_out<=8'b00010001;
        13'd1482: m_out<=8'b00010010;
        13'd1483: m_out<=8'b00001010;
        13'd1484: m_out<=8'b00000001;
        13'd1485: m_out<=8'b00101000;
        13'd1486: m_out<=8'b00000110;
        13'd1487: m_out<=8'b00000001;
        13'd1488: m_out<=8'b11110000;
        13'd1489: m_out<=8'b00000111;
        13'd1490: m_out<=8'b00010011;
        13'd1491: m_out<=8'b11010101;
        13'd1492: m_out<=8'b00100001;
        13'd1493: m_out<=8'b00000111;
        13'd1494: m_out<=8'b11100000;
        13'd1495: m_out<=8'b00100000;
        13'd1496: m_out<=8'b00000111;
        13'd1497: m_out<=8'b00010100;
        13'd1498: m_out<=8'b11111100;
        13'd1499: m_out<=8'b11110111;
        13'd1500: m_out<=8'b11110110;
        13'd1501: m_out<=8'b00011011;
        13'd1502: m_out<=8'b00000111;
        13'd1503: m_out<=8'b11011110;
        13'd1504: m_out<=8'b00001110;
        13'd1505: m_out<=8'b11100100;
        13'd1506: m_out<=8'b00011000;
        13'd1507: m_out<=8'b00000111;
        13'd1508: m_out<=8'b11100111;
        13'd1509: m_out<=8'b11110011;
        13'd1510: m_out<=8'b11011100;
        13'd1511: m_out<=8'b00010010;
        13'd1512: m_out<=8'b00010101;
        13'd1513: m_out<=8'b00001111;
        13'd1514: m_out<=8'b00100001;
        13'd1515: m_out<=8'b00100001;
        13'd1516: m_out<=8'b00001010;
        13'd1517: m_out<=8'b11011110;
        13'd1518: m_out<=8'b11111110;
        13'd1519: m_out<=8'b00000011;
        13'd1520: m_out<=8'b00000000;
        13'd1521: m_out<=8'b11011110;
        13'd1522: m_out<=8'b11101011;
        13'd1523: m_out<=8'b11111101;
        13'd1524: m_out<=8'b00100000;
        13'd1525: m_out<=8'b00010100;
        13'd1526: m_out<=8'b00011010;
        13'd1527: m_out<=8'b11111000;
        13'd1528: m_out<=8'b11110101;
        13'd1529: m_out<=8'b00011010;
        13'd1530: m_out<=8'b00000001;
        13'd1531: m_out<=8'b11101101;
        13'd1532: m_out<=8'b11110010;
        13'd1533: m_out<=8'b11110010;
        13'd1534: m_out<=8'b00100001;
        13'd1535: m_out<=8'b00001101;
        13'd1536: m_out<=8'b00000000;
        13'd1537: m_out<=8'b00000011;
        13'd1538: m_out<=8'b00000111;
        13'd1539: m_out<=8'b00011111;
        13'd1540: m_out<=8'b00001011;
        13'd1541: m_out<=8'b11100101;
        13'd1542: m_out<=8'b11100111;
        13'd1543: m_out<=8'b00001101;
        13'd1544: m_out<=8'b00001000;
        13'd1545: m_out<=8'b11111010;
        13'd1546: m_out<=8'b11010100;
        13'd1547: m_out<=8'b00100100;
        13'd1548: m_out<=8'b11101110;
        13'd1549: m_out<=8'b00101101;
        13'd1550: m_out<=8'b00000011;
        13'd1551: m_out<=8'b11110011;
        13'd1552: m_out<=8'b11101100;
        13'd1553: m_out<=8'b11100110;
        13'd1554: m_out<=8'b11011010;
        13'd1555: m_out<=8'b11010110;
        13'd1556: m_out<=8'b00010001;
        13'd1557: m_out<=8'b11111000;
        13'd1558: m_out<=8'b00001101;
        13'd1559: m_out<=8'b11100111;
        13'd1560: m_out<=8'b00001010;
        13'd1561: m_out<=8'b11111100;
        13'd1562: m_out<=8'b00000101;
        13'd1563: m_out<=8'b00111110;
        13'd1564: m_out<=8'b00010011;
        13'd1565: m_out<=8'b11101010;
        13'd1566: m_out<=8'b11110110;
        13'd1567: m_out<=8'b11111001;
        13'd1568: m_out<=8'b11100011;
        13'd1569: m_out<=8'b11101101;
        13'd1570: m_out<=8'b11101100;
        13'd1571: m_out<=8'b11110101;
        13'd1572: m_out<=8'b00000001;
        13'd1573: m_out<=8'b00001100;
        13'd1574: m_out<=8'b11100111;
        13'd1575: m_out<=8'b00001110;
        13'd1576: m_out<=8'b00000110;
        13'd1577: m_out<=8'b00010000;
        13'd1578: m_out<=8'b00011101;
        13'd1579: m_out<=8'b11100101;
        13'd1580: m_out<=8'b00110111;
        13'd1581: m_out<=8'b11011000;
        13'd1582: m_out<=8'b00011001;
        13'd1583: m_out<=8'b11011010;
        13'd1584: m_out<=8'b00011011;
        13'd1585: m_out<=8'b00001001;
        13'd1586: m_out<=8'b00110111;
        13'd1587: m_out<=8'b11110110;
        13'd1588: m_out<=8'b11010001;
        13'd1589: m_out<=8'b00000100;
        13'd1590: m_out<=8'b11110100;
        13'd1591: m_out<=8'b00001100;
        13'd1592: m_out<=8'b11110010;
        13'd1593: m_out<=8'b11110000;
        13'd1594: m_out<=8'b11100111;
        13'd1595: m_out<=8'b11110100;
        13'd1596: m_out<=8'b11100110;
        13'd1597: m_out<=8'b00010011;
        13'd1598: m_out<=8'b11111100;
        13'd1599: m_out<=8'b11111000;
        13'd1600: m_out<=8'b11101100;
        13'd1601: m_out<=8'b00100000;
        13'd1602: m_out<=8'b00011011;
        13'd1603: m_out<=8'b00010001;
        13'd1604: m_out<=8'b11110101;
        13'd1605: m_out<=8'b00011001;
        13'd1606: m_out<=8'b11011101;
        13'd1607: m_out<=8'b00010101;
        13'd1608: m_out<=8'b11100111;
        13'd1609: m_out<=8'b00000001;
        13'd1610: m_out<=8'b11101111;
        13'd1611: m_out<=8'b11011111;
        13'd1612: m_out<=8'b00010000;
        13'd1613: m_out<=8'b11010011;
        13'd1614: m_out<=8'b11110111;
        13'd1615: m_out<=8'b11111110;
        13'd1616: m_out<=8'b00111000;
        13'd1617: m_out<=8'b00000000;
        13'd1618: m_out<=8'b00001110;
        13'd1619: m_out<=8'b11110001;
        13'd1620: m_out<=8'b11011110;
        13'd1621: m_out<=8'b00000011;
        13'd1622: m_out<=8'b11100111;
        13'd1623: m_out<=8'b11111110;
        13'd1624: m_out<=8'b11110011;
        13'd1625: m_out<=8'b00001111;
        13'd1626: m_out<=8'b00001101;
        13'd1627: m_out<=8'b00100100;
        13'd1628: m_out<=8'b11110001;
        13'd1629: m_out<=8'b00100100;
        13'd1630: m_out<=8'b11111101;
        13'd1631: m_out<=8'b11111100;
        13'd1632: m_out<=8'b00010110;
        13'd1633: m_out<=8'b11100010;
        13'd1634: m_out<=8'b00010111;
        13'd1635: m_out<=8'b11001111;
        13'd1636: m_out<=8'b11011000;
        13'd1637: m_out<=8'b11110100;
        13'd1638: m_out<=8'b00001100;
        13'd1639: m_out<=8'b00001100;
        13'd1640: m_out<=8'b11111001;
        13'd1641: m_out<=8'b00001001;
        13'd1642: m_out<=8'b00001010;
        13'd1643: m_out<=8'b11101110;
        13'd1644: m_out<=8'b00000010;
        13'd1645: m_out<=8'b00001100;
        13'd1646: m_out<=8'b00101001;
        13'd1647: m_out<=8'b11100111;
        13'd1648: m_out<=8'b00001001;
        13'd1649: m_out<=8'b00001010;
        13'd1650: m_out<=8'b00011100;
        13'd1651: m_out<=8'b00011100;
        13'd1652: m_out<=8'b00001110;
        13'd1653: m_out<=8'b11101100;
        13'd1654: m_out<=8'b00000110;
        13'd1655: m_out<=8'b11111010;
        13'd1656: m_out<=8'b11001010;
        13'd1657: m_out<=8'b11000100;
        13'd1658: m_out<=8'b00010011;
        13'd1659: m_out<=8'b00001100;
        13'd1660: m_out<=8'b11010111;
        13'd1661: m_out<=8'b10111111;
        13'd1662: m_out<=8'b11101000;
        13'd1663: m_out<=8'b11011000;
        13'd1664: m_out<=8'b00010101;
        13'd1665: m_out<=8'b00001100;
        13'd1666: m_out<=8'b11100110;
        13'd1667: m_out<=8'b11110100;
        13'd1668: m_out<=8'b00000110;
        13'd1669: m_out<=8'b11010000;
        13'd1670: m_out<=8'b00111000;
        13'd1671: m_out<=8'b00100110;
        13'd1672: m_out<=8'b00001001;
        13'd1673: m_out<=8'b11010010;
        13'd1674: m_out<=8'b00011001;
        13'd1675: m_out<=8'b11111011;
        13'd1676: m_out<=8'b11110101;
        13'd1677: m_out<=8'b00001100;
        13'd1678: m_out<=8'b11110001;
        13'd1679: m_out<=8'b00100000;
        13'd1680: m_out<=8'b11011110;
        13'd1681: m_out<=8'b11110100;
        13'd1682: m_out<=8'b11100000;
        13'd1683: m_out<=8'b00110000;
        13'd1684: m_out<=8'b00000010;
        13'd1685: m_out<=8'b00110001;
        13'd1686: m_out<=8'b11110001;
        13'd1687: m_out<=8'b11110011;
        13'd1688: m_out<=8'b11010011;
        13'd1689: m_out<=8'b11010101;
        13'd1690: m_out<=8'b11110010;
        13'd1691: m_out<=8'b00000011;
        13'd1692: m_out<=8'b00000100;
        13'd1693: m_out<=8'b11100011;
        13'd1694: m_out<=8'b11100111;
        13'd1695: m_out<=8'b00011101;
        13'd1696: m_out<=8'b00000101;
        13'd1697: m_out<=8'b00111011;
        13'd1698: m_out<=8'b00100101;
        13'd1699: m_out<=8'b11010000;
        13'd1700: m_out<=8'b00001001;
        13'd1701: m_out<=8'b11100110;
        13'd1702: m_out<=8'b11000110;
        13'd1703: m_out<=8'b11111101;
        13'd1704: m_out<=8'b11111010;
        13'd1705: m_out<=8'b11111100;
        13'd1706: m_out<=8'b00010111;
        13'd1707: m_out<=8'b11111101;
        13'd1708: m_out<=8'b00000100;
        13'd1709: m_out<=8'b11110000;
        13'd1710: m_out<=8'b00000001;
        13'd1711: m_out<=8'b00000000;
        13'd1712: m_out<=8'b11110001;
        13'd1713: m_out<=8'b00000101;
        13'd1714: m_out<=8'b00000101;
        13'd1715: m_out<=8'b00001001;
        13'd1716: m_out<=8'b11100100;
        13'd1717: m_out<=8'b00010001;
        13'd1718: m_out<=8'b11110111;
        13'd1719: m_out<=8'b00001100;
        13'd1720: m_out<=8'b11101000;
        13'd1721: m_out<=8'b11110101;
        13'd1722: m_out<=8'b11010111;
        13'd1723: m_out<=8'b11110100;
        13'd1724: m_out<=8'b00100001;
        13'd1725: m_out<=8'b11000101;
        13'd1726: m_out<=8'b11111111;
        13'd1727: m_out<=8'b11110100;
        13'd1728: m_out<=8'b11111000;
        13'd1729: m_out<=8'b00101011;
        13'd1730: m_out<=8'b11110111;
        13'd1731: m_out<=8'b11011111;
        13'd1732: m_out<=8'b11110110;
        13'd1733: m_out<=8'b00000111;
        13'd1734: m_out<=8'b00001010;
        13'd1735: m_out<=8'b00011110;
        13'd1736: m_out<=8'b11111101;
        13'd1737: m_out<=8'b00110010;
        13'd1738: m_out<=8'b11100110;
        13'd1739: m_out<=8'b00000100;
        13'd1740: m_out<=8'b00000101;
        13'd1741: m_out<=8'b11111010;
        13'd1742: m_out<=8'b00010010;
        13'd1743: m_out<=8'b11000110;
        13'd1744: m_out<=8'b11111000;
        13'd1745: m_out<=8'b11101010;
        13'd1746: m_out<=8'b11110100;
        13'd1747: m_out<=8'b11101101;
        13'd1748: m_out<=8'b11100001;
        13'd1749: m_out<=8'b11101101;
        13'd1750: m_out<=8'b00000101;
        13'd1751: m_out<=8'b11110110;
        13'd1752: m_out<=8'b11011001;
        13'd1753: m_out<=8'b00001000;
        13'd1754: m_out<=8'b11111111;
        13'd1755: m_out<=8'b00001111;
        13'd1756: m_out<=8'b11101001;
        13'd1757: m_out<=8'b11111110;
        13'd1758: m_out<=8'b11111110;
        13'd1759: m_out<=8'b11110000;
        13'd1760: m_out<=8'b00011100;
        13'd1761: m_out<=8'b11110100;
        13'd1762: m_out<=8'b00010111;
        13'd1763: m_out<=8'b00000001;
        13'd1764: m_out<=8'b00000101;
        13'd1765: m_out<=8'b11010011;
        13'd1766: m_out<=8'b11100111;
        13'd1767: m_out<=8'b00000010;
        13'd1768: m_out<=8'b00011010;
        13'd1769: m_out<=8'b00000110;
        13'd1770: m_out<=8'b00000110;
        13'd1771: m_out<=8'b00011011;
        13'd1772: m_out<=8'b00000010;
        13'd1773: m_out<=8'b00111110;
        13'd1774: m_out<=8'b11110011;
        13'd1775: m_out<=8'b11101100;
        13'd1776: m_out<=8'b00000100;
        13'd1777: m_out<=8'b00101011;
        13'd1778: m_out<=8'b11101101;
        13'd1779: m_out<=8'b11110101;
        13'd1780: m_out<=8'b00101101;
        13'd1781: m_out<=8'b00100010;
        13'd1782: m_out<=8'b00101100;
        13'd1783: m_out<=8'b11011100;
        13'd1784: m_out<=8'b00001001;
        13'd1785: m_out<=8'b11100001;
        13'd1786: m_out<=8'b11100101;
        13'd1787: m_out<=8'b11101011;
        13'd1788: m_out<=8'b11110111;
        13'd1789: m_out<=8'b11101111;
        13'd1790: m_out<=8'b11011011;
        13'd1791: m_out<=8'b00000101;
        13'd1792: m_out<=8'b11111101;
        13'd1793: m_out<=8'b00000010;
        13'd1794: m_out<=8'b00011100;
        13'd1795: m_out<=8'b11110111;
        13'd1796: m_out<=8'b10111011;
        13'd1797: m_out<=8'b00000010;
        13'd1798: m_out<=8'b00010010;
        13'd1799: m_out<=8'b00100100;
        13'd1800: m_out<=8'b00001100;
        13'd1801: m_out<=8'b11110110;
        13'd1802: m_out<=8'b00111010;
        13'd1803: m_out<=8'b11111011;
        13'd1804: m_out<=8'b00001110;
        13'd1805: m_out<=8'b11101101;
        13'd1806: m_out<=8'b00000111;
        13'd1807: m_out<=8'b11111100;
        13'd1808: m_out<=8'b00001001;
        13'd1809: m_out<=8'b11010010;
        13'd1810: m_out<=8'b00010101;
        13'd1811: m_out<=8'b11110100;
        13'd1812: m_out<=8'b00000100;
        13'd1813: m_out<=8'b00001110;
        13'd1814: m_out<=8'b00001010;
        13'd1815: m_out<=8'b00001001;
        13'd1816: m_out<=8'b11110111;
        13'd1817: m_out<=8'b11100000;
        13'd1818: m_out<=8'b11101011;
        13'd1819: m_out<=8'b11111110;
        13'd1820: m_out<=8'b00001011;
        13'd1821: m_out<=8'b11110111;
        13'd1822: m_out<=8'b11110000;
        13'd1823: m_out<=8'b00000011;
        13'd1824: m_out<=8'b00010110;
        13'd1825: m_out<=8'b00010111;
        13'd1826: m_out<=8'b11110010;
        13'd1827: m_out<=8'b00001111;
        13'd1828: m_out<=8'b11100101;
        13'd1829: m_out<=8'b11101110;
        13'd1830: m_out<=8'b00011010;
        13'd1831: m_out<=8'b11000101;
        13'd1832: m_out<=8'b11100100;
        13'd1833: m_out<=8'b00100001;
        13'd1834: m_out<=8'b00001001;
        13'd1835: m_out<=8'b11100101;
        13'd1836: m_out<=8'b11110101;
        13'd1837: m_out<=8'b11110111;
        13'd1838: m_out<=8'b00011111;
        13'd1839: m_out<=8'b11111110;
        13'd1840: m_out<=8'b00110101;
        13'd1841: m_out<=8'b00100011;
        13'd1842: m_out<=8'b11010100;
        13'd1843: m_out<=8'b00101001;
        13'd1844: m_out<=8'b00000110;
        13'd1845: m_out<=8'b00001000;
        13'd1846: m_out<=8'b00101000;
        13'd1847: m_out<=8'b00000010;
        13'd1848: m_out<=8'b00100110;
        13'd1849: m_out<=8'b00011011;
        13'd1850: m_out<=8'b00000101;
        13'd1851: m_out<=8'b11101001;
        13'd1852: m_out<=8'b11111101;
        13'd1853: m_out<=8'b11011011;
        13'd1854: m_out<=8'b00001011;
        13'd1855: m_out<=8'b00000100;
        13'd1856: m_out<=8'b11100111;
        13'd1857: m_out<=8'b00000000;
        13'd1858: m_out<=8'b00100111;
        13'd1859: m_out<=8'b00011010;
        13'd1860: m_out<=8'b11011010;
        13'd1861: m_out<=8'b11111000;
        13'd1862: m_out<=8'b00001011;
        13'd1863: m_out<=8'b00001100;
        13'd1864: m_out<=8'b11100000;
        13'd1865: m_out<=8'b00001011;
        13'd1866: m_out<=8'b00001110;
        13'd1867: m_out<=8'b00000001;
        13'd1868: m_out<=8'b00101011;
        13'd1869: m_out<=8'b11110110;
        13'd1870: m_out<=8'b11111111;
        13'd1871: m_out<=8'b00000010;
        13'd1872: m_out<=8'b00011000;
        13'd1873: m_out<=8'b11101100;
        13'd1874: m_out<=8'b00010111;
        13'd1875: m_out<=8'b11110110;
        13'd1876: m_out<=8'b00001100;
        13'd1877: m_out<=8'b11101100;
        13'd1878: m_out<=8'b00001010;
        13'd1879: m_out<=8'b00010111;
        13'd1880: m_out<=8'b11011110;
        13'd1881: m_out<=8'b11101110;
        13'd1882: m_out<=8'b11110111;
        13'd1883: m_out<=8'b11110110;
        13'd1884: m_out<=8'b11100101;
        13'd1885: m_out<=8'b00000010;
        13'd1886: m_out<=8'b11111011;
        13'd1887: m_out<=8'b00100010;
        13'd1888: m_out<=8'b11111110;
        13'd1889: m_out<=8'b00101101;
        13'd1890: m_out<=8'b11100011;
        13'd1891: m_out<=8'b11000011;
        13'd1892: m_out<=8'b11111000;
        13'd1893: m_out<=8'b00011001;
        13'd1894: m_out<=8'b11110110;
        13'd1895: m_out<=8'b11111111;
        13'd1896: m_out<=8'b11101011;
        13'd1897: m_out<=8'b11110111;
        13'd1898: m_out<=8'b11101010;
        13'd1899: m_out<=8'b11111101;
        13'd1900: m_out<=8'b11101100;
        13'd1901: m_out<=8'b11101100;
        13'd1902: m_out<=8'b00010000;
        13'd1903: m_out<=8'b11110000;
        13'd1904: m_out<=8'b00011100;
        13'd1905: m_out<=8'b00001111;
        13'd1906: m_out<=8'b00011111;
        13'd1907: m_out<=8'b11011101;
        13'd1908: m_out<=8'b11110000;
        13'd1909: m_out<=8'b00000010;
        13'd1910: m_out<=8'b11000111;
        13'd1911: m_out<=8'b11111111;
        13'd1912: m_out<=8'b11110000;
        13'd1913: m_out<=8'b11100101;
        13'd1914: m_out<=8'b00000000;
        13'd1915: m_out<=8'b11110110;
        13'd1916: m_out<=8'b00100101;
        13'd1917: m_out<=8'b00000100;
        13'd1918: m_out<=8'b00000101;
        13'd1919: m_out<=8'b11110010;
        13'd1920: m_out<=8'b11111001;
        13'd1921: m_out<=8'b11110010;
        13'd1922: m_out<=8'b11101001;
        13'd1923: m_out<=8'b11110110;
        13'd1924: m_out<=8'b00001110;
        13'd1925: m_out<=8'b11011110;
        13'd1926: m_out<=8'b00000111;
        13'd1927: m_out<=8'b11101101;
        13'd1928: m_out<=8'b00110100;
        13'd1929: m_out<=8'b00001011;
        13'd1930: m_out<=8'b00000110;
        13'd1931: m_out<=8'b00011011;
        13'd1932: m_out<=8'b11110111;
        13'd1933: m_out<=8'b11000111;
        13'd1934: m_out<=8'b11100101;
        13'd1935: m_out<=8'b00011001;
        13'd1936: m_out<=8'b00010101;
        13'd1937: m_out<=8'b00000000;
        13'd1938: m_out<=8'b11111100;
        13'd1939: m_out<=8'b11100100;
        13'd1940: m_out<=8'b11110101;
        13'd1941: m_out<=8'b11011110;
        13'd1942: m_out<=8'b11101011;
        13'd1943: m_out<=8'b00010001;
        13'd1944: m_out<=8'b11101100;
        13'd1945: m_out<=8'b00001010;
        13'd1946: m_out<=8'b11110011;
        13'd1947: m_out<=8'b11111011;
        13'd1948: m_out<=8'b00010110;
        13'd1949: m_out<=8'b00001001;
        13'd1950: m_out<=8'b00100111;
        13'd1951: m_out<=8'b11100100;
        13'd1952: m_out<=8'b00000111;
        13'd1953: m_out<=8'b00000101;
        13'd1954: m_out<=8'b11101111;
        13'd1955: m_out<=8'b11100001;
        13'd1956: m_out<=8'b11001100;
        13'd1957: m_out<=8'b00110111;
        13'd1958: m_out<=8'b11101100;
        13'd1959: m_out<=8'b00010000;
        13'd1960: m_out<=8'b00010001;
        13'd1961: m_out<=8'b11111011;
        13'd1962: m_out<=8'b00010010;
        13'd1963: m_out<=8'b00000100;
        13'd1964: m_out<=8'b11110011;
        13'd1965: m_out<=8'b00010101;
        13'd1966: m_out<=8'b00010110;
        13'd1967: m_out<=8'b11100101;
        13'd1968: m_out<=8'b10111011;
        13'd1969: m_out<=8'b11111110;
        13'd1970: m_out<=8'b11111100;
        13'd1971: m_out<=8'b00010011;
        13'd1972: m_out<=8'b11110110;
        13'd1973: m_out<=8'b00000000;
        13'd1974: m_out<=8'b00000110;
        13'd1975: m_out<=8'b11101010;
        13'd1976: m_out<=8'b00011001;
        13'd1977: m_out<=8'b00100001;
        13'd1978: m_out<=8'b00001111;
        13'd1979: m_out<=8'b00110101;
        13'd1980: m_out<=8'b11111001;
        13'd1981: m_out<=8'b11110001;
        13'd1982: m_out<=8'b00101000;
        13'd1983: m_out<=8'b00010010;
        13'd1984: m_out<=8'b11100001;
        13'd1985: m_out<=8'b11010010;
        13'd1986: m_out<=8'b11110111;
        13'd1987: m_out<=8'b00001110;
        13'd1988: m_out<=8'b11100010;
        13'd1989: m_out<=8'b11101010;
        13'd1990: m_out<=8'b00001000;
        13'd1991: m_out<=8'b11011011;
        13'd1992: m_out<=8'b00000100;
        13'd1993: m_out<=8'b11110011;
        13'd1994: m_out<=8'b11110110;
        13'd1995: m_out<=8'b11010110;
        13'd1996: m_out<=8'b00001100;
        13'd1997: m_out<=8'b00101001;
        13'd1998: m_out<=8'b00001011;
        13'd1999: m_out<=8'b00001101;
        13'd2000: m_out<=8'b00010111;
        13'd2001: m_out<=8'b00000110;
        13'd2002: m_out<=8'b10111010;
        13'd2003: m_out<=8'b00001101;
        13'd2004: m_out<=8'b00100000;
        13'd2005: m_out<=8'b00001101;
        13'd2006: m_out<=8'b11010010;
        13'd2007: m_out<=8'b00000101;
        13'd2008: m_out<=8'b11101110;
        13'd2009: m_out<=8'b00010001;
        13'd2010: m_out<=8'b11111000;
        13'd2011: m_out<=8'b00001010;
        13'd2012: m_out<=8'b11111010;
        13'd2013: m_out<=8'b00000100;
        13'd2014: m_out<=8'b11110101;
        13'd2015: m_out<=8'b00111110;
        13'd2016: m_out<=8'b00010000;
        13'd2017: m_out<=8'b11100010;
        13'd2018: m_out<=8'b00001001;
        13'd2019: m_out<=8'b00010000;
        13'd2020: m_out<=8'b11110010;
        13'd2021: m_out<=8'b11110110;
        13'd2022: m_out<=8'b11111110;
        13'd2023: m_out<=8'b00001100;
        13'd2024: m_out<=8'b00001100;
        13'd2025: m_out<=8'b10111010;
        13'd2026: m_out<=8'b11110001;
        13'd2027: m_out<=8'b11100101;
        13'd2028: m_out<=8'b11110010;
        13'd2029: m_out<=8'b11101011;
        13'd2030: m_out<=8'b11111110;
        13'd2031: m_out<=8'b00100000;
        13'd2032: m_out<=8'b11101110;
        13'd2033: m_out<=8'b11011111;
        13'd2034: m_out<=8'b00001111;
        13'd2035: m_out<=8'b11110000;
        13'd2036: m_out<=8'b00000011;
        13'd2037: m_out<=8'b11001010;
        13'd2038: m_out<=8'b00111111;
        13'd2039: m_out<=8'b11110101;
        13'd2040: m_out<=8'b00110010;
        13'd2041: m_out<=8'b11101011;
        13'd2042: m_out<=8'b11100101;
        13'd2043: m_out<=8'b00010100;
        13'd2044: m_out<=8'b11101111;
        13'd2045: m_out<=8'b00001110;
        13'd2046: m_out<=8'b00001111;
        13'd2047: m_out<=8'b11001111;
        13'd2048: m_out<=8'b00111001;
        13'd2049: m_out<=8'b11101100;
        13'd2050: m_out<=8'b11111010;
        13'd2051: m_out<=8'b11111011;
        13'd2052: m_out<=8'b00010111;
        13'd2053: m_out<=8'b11011100;
        13'd2054: m_out<=8'b00000011;
        13'd2055: m_out<=8'b00010001;
        13'd2056: m_out<=8'b00000111;
        13'd2057: m_out<=8'b00011110;
        13'd2058: m_out<=8'b11111100;
        13'd2059: m_out<=8'b11110011;
        13'd2060: m_out<=8'b00100010;
        13'd2061: m_out<=8'b11111110;
        13'd2062: m_out<=8'b11111110;
        13'd2063: m_out<=8'b11010110;
        13'd2064: m_out<=8'b00011010;
        13'd2065: m_out<=8'b11001010;
        13'd2066: m_out<=8'b00010001;
        13'd2067: m_out<=8'b11010010;
        13'd2068: m_out<=8'b11110111;
        13'd2069: m_out<=8'b11001110;
        13'd2070: m_out<=8'b00011001;
        13'd2071: m_out<=8'b00001101;
        13'd2072: m_out<=8'b11101000;
        13'd2073: m_out<=8'b11000111;
        13'd2074: m_out<=8'b00000001;
        13'd2075: m_out<=8'b11110100;
        13'd2076: m_out<=8'b11001001;
        13'd2077: m_out<=8'b11100100;
        13'd2078: m_out<=8'b00010001;
        13'd2079: m_out<=8'b00000001;
        13'd2080: m_out<=8'b11101001;
        13'd2081: m_out<=8'b00110011;
        13'd2082: m_out<=8'b00001011;
        13'd2083: m_out<=8'b00000000;
        13'd2084: m_out<=8'b00000110;
        13'd2085: m_out<=8'b00000011;
        13'd2086: m_out<=8'b00001111;
        13'd2087: m_out<=8'b11110110;
        13'd2088: m_out<=8'b11011111;
        13'd2089: m_out<=8'b11001101;
        13'd2090: m_out<=8'b00000110;
        13'd2091: m_out<=8'b11111111;
        13'd2092: m_out<=8'b00001001;
        13'd2093: m_out<=8'b11110111;
        13'd2094: m_out<=8'b11111111;
        13'd2095: m_out<=8'b11101101;
        13'd2096: m_out<=8'b00001100;
        13'd2097: m_out<=8'b00101010;
        13'd2098: m_out<=8'b00010101;
        13'd2099: m_out<=8'b00011010;
        13'd2100: m_out<=8'b00110100;
        13'd2101: m_out<=8'b11111101;
        13'd2102: m_out<=8'b11111010;
        13'd2103: m_out<=8'b00000100;
        13'd2104: m_out<=8'b00000011;
        13'd2105: m_out<=8'b11110101;
        13'd2106: m_out<=8'b11110101;
        13'd2107: m_out<=8'b11110101;
        13'd2108: m_out<=8'b11100100;
        13'd2109: m_out<=8'b00000101;
        13'd2110: m_out<=8'b11100101;
        13'd2111: m_out<=8'b00000000;
        13'd2112: m_out<=8'b00110101;
        13'd2113: m_out<=8'b00010011;
        13'd2114: m_out<=8'b11110010;
        13'd2115: m_out<=8'b11011100;
        13'd2116: m_out<=8'b00000010;
        13'd2117: m_out<=8'b11110101;
        13'd2118: m_out<=8'b11011011;
        13'd2119: m_out<=8'b00011101;
        13'd2120: m_out<=8'b11111101;
        13'd2121: m_out<=8'b11110011;
        13'd2122: m_out<=8'b11101111;
        13'd2123: m_out<=8'b00001000;
        13'd2124: m_out<=8'b00010110;
        13'd2125: m_out<=8'b00011011;
        13'd2126: m_out<=8'b11101110;
        13'd2127: m_out<=8'b11110010;
        13'd2128: m_out<=8'b00011011;
        13'd2129: m_out<=8'b11101111;
        13'd2130: m_out<=8'b00101101;
        13'd2131: m_out<=8'b00011010;
        13'd2132: m_out<=8'b11100101;
        13'd2133: m_out<=8'b00001100;
        13'd2134: m_out<=8'b00000110;
        13'd2135: m_out<=8'b11110100;
        13'd2136: m_out<=8'b00011111;
        13'd2137: m_out<=8'b00011101;
        13'd2138: m_out<=8'b00001111;
        13'd2139: m_out<=8'b11110111;
        13'd2140: m_out<=8'b11111100;
        13'd2141: m_out<=8'b00000100;
        13'd2142: m_out<=8'b11110110;
        13'd2143: m_out<=8'b00001000;
        13'd2144: m_out<=8'b01000001;
        13'd2145: m_out<=8'b00001010;
        13'd2146: m_out<=8'b11100110;
        13'd2147: m_out<=8'b11110111;
        13'd2148: m_out<=8'b00001101;
        13'd2149: m_out<=8'b00011000;
        13'd2150: m_out<=8'b00000101;
        13'd2151: m_out<=8'b00010010;
        13'd2152: m_out<=8'b11111111;
        13'd2153: m_out<=8'b00010011;
        13'd2154: m_out<=8'b11110111;
        13'd2155: m_out<=8'b11110100;
        13'd2156: m_out<=8'b00011110;
        13'd2157: m_out<=8'b00010011;
        13'd2158: m_out<=8'b11111000;
        13'd2159: m_out<=8'b11100010;
        13'd2160: m_out<=8'b11101101;
        13'd2161: m_out<=8'b11100101;
        13'd2162: m_out<=8'b00100000;
        13'd2163: m_out<=8'b11011010;
        13'd2164: m_out<=8'b00010011;
        13'd2165: m_out<=8'b11010101;
        13'd2166: m_out<=8'b11111100;
        13'd2167: m_out<=8'b00101111;
        13'd2168: m_out<=8'b00100100;
        13'd2169: m_out<=8'b11101110;
        13'd2170: m_out<=8'b00010001;
        13'd2171: m_out<=8'b11100100;
        13'd2172: m_out<=8'b00010000;
        13'd2173: m_out<=8'b11001111;
        13'd2174: m_out<=8'b11100111;
        13'd2175: m_out<=8'b11101111;
        13'd2176: m_out<=8'b00000110;
        13'd2177: m_out<=8'b11100011;
        13'd2178: m_out<=8'b11111110;
        13'd2179: m_out<=8'b11110010;
        13'd2180: m_out<=8'b00010011;
        13'd2181: m_out<=8'b11101100;
        13'd2182: m_out<=8'b00010010;
        13'd2183: m_out<=8'b11011110;
        13'd2184: m_out<=8'b11101111;
        13'd2185: m_out<=8'b00001001;
        13'd2186: m_out<=8'b00010111;
        13'd2187: m_out<=8'b00010010;
        13'd2188: m_out<=8'b11111101;
        13'd2189: m_out<=8'b00011000;
        13'd2190: m_out<=8'b00000111;
        13'd2191: m_out<=8'b11010111;
        13'd2192: m_out<=8'b11011111;
        13'd2193: m_out<=8'b00000001;
        13'd2194: m_out<=8'b00000010;
        13'd2195: m_out<=8'b11100010;
        13'd2196: m_out<=8'b00000000;
        13'd2197: m_out<=8'b00001011;
        13'd2198: m_out<=8'b11100011;
        13'd2199: m_out<=8'b00100001;
        13'd2200: m_out<=8'b11111010;
        13'd2201: m_out<=8'b00100000;
        13'd2202: m_out<=8'b11010010;
        13'd2203: m_out<=8'b00001000;
        13'd2204: m_out<=8'b11011100;
        13'd2205: m_out<=8'b00010100;
        13'd2206: m_out<=8'b00011111;
        13'd2207: m_out<=8'b11101000;
        13'd2208: m_out<=8'b11110001;
        13'd2209: m_out<=8'b11100101;
        13'd2210: m_out<=8'b11111000;
        13'd2211: m_out<=8'b11011001;
        13'd2212: m_out<=8'b11111001;
        13'd2213: m_out<=8'b00000100;
        13'd2214: m_out<=8'b11110111;
        13'd2215: m_out<=8'b00001001;
        13'd2216: m_out<=8'b00001001;
        13'd2217: m_out<=8'b11010101;
        13'd2218: m_out<=8'b00011110;
        13'd2219: m_out<=8'b11111010;
        13'd2220: m_out<=8'b11100101;
        13'd2221: m_out<=8'b11101001;
        13'd2222: m_out<=8'b00000110;
        13'd2223: m_out<=8'b11110011;
        13'd2224: m_out<=8'b11111010;
        13'd2225: m_out<=8'b11101101;
        13'd2226: m_out<=8'b11011001;
        13'd2227: m_out<=8'b00010110;
        13'd2228: m_out<=8'b11110100;
        13'd2229: m_out<=8'b00100101;
        13'd2230: m_out<=8'b11110111;
        13'd2231: m_out<=8'b00011101;
        13'd2232: m_out<=8'b00011110;
        13'd2233: m_out<=8'b00010100;
        13'd2234: m_out<=8'b00011100;
        13'd2235: m_out<=8'b00010001;
        13'd2236: m_out<=8'b00100101;
        13'd2237: m_out<=8'b11110100;
        13'd2238: m_out<=8'b00000111;
        13'd2239: m_out<=8'b00101101;
        13'd2240: m_out<=8'b00011001;
        13'd2241: m_out<=8'b11000111;
        13'd2242: m_out<=8'b11100000;
        13'd2243: m_out<=8'b11111000;
        13'd2244: m_out<=8'b11101010;
        13'd2245: m_out<=8'b00100110;
        13'd2246: m_out<=8'b00101000;
        13'd2247: m_out<=8'b11001001;
        13'd2248: m_out<=8'b11000101;
        13'd2249: m_out<=8'b00001001;
        13'd2250: m_out<=8'b11110100;
        13'd2251: m_out<=8'b00001101;
        13'd2252: m_out<=8'b00010001;
        13'd2253: m_out<=8'b00001111;
        13'd2254: m_out<=8'b00000001;
        13'd2255: m_out<=8'b11110100;
        13'd2256: m_out<=8'b11101101;
        13'd2257: m_out<=8'b11010001;
        13'd2258: m_out<=8'b11100001;
        13'd2259: m_out<=8'b00001000;
        13'd2260: m_out<=8'b00100101;
        13'd2261: m_out<=8'b00100101;
        13'd2262: m_out<=8'b00011100;
        13'd2263: m_out<=8'b11110000;
        13'd2264: m_out<=8'b11011100;
        13'd2265: m_out<=8'b11001110;
        13'd2266: m_out<=8'b00111101;
        13'd2267: m_out<=8'b11101100;
        13'd2268: m_out<=8'b00111010;
        13'd2269: m_out<=8'b00110011;
        13'd2270: m_out<=8'b00000011;
        13'd2271: m_out<=8'b11011011;
        13'd2272: m_out<=8'b11010011;
        13'd2273: m_out<=8'b00000101;
        13'd2274: m_out<=8'b11011110;
        13'd2275: m_out<=8'b11011001;
        13'd2276: m_out<=8'b00100001;
        13'd2277: m_out<=8'b11110011;
        13'd2278: m_out<=8'b00100000;
        13'd2279: m_out<=8'b11111000;
        13'd2280: m_out<=8'b00010100;
        13'd2281: m_out<=8'b11110010;
        13'd2282: m_out<=8'b11111101;
        13'd2283: m_out<=8'b00101111;
        13'd2284: m_out<=8'b11111101;
        13'd2285: m_out<=8'b11111111;
        13'd2286: m_out<=8'b00011100;
        13'd2287: m_out<=8'b00000001;
        13'd2288: m_out<=8'b00110110;
        13'd2289: m_out<=8'b11110110;
        13'd2290: m_out<=8'b00011111;
        13'd2291: m_out<=8'b00001111;
        13'd2292: m_out<=8'b11000110;
        13'd2293: m_out<=8'b00001011;
        13'd2294: m_out<=8'b00001111;
        13'd2295: m_out<=8'b00001111;
        13'd2296: m_out<=8'b11110000;
        13'd2297: m_out<=8'b11011001;
        13'd2298: m_out<=8'b00001001;
        13'd2299: m_out<=8'b00000101;
        13'd2300: m_out<=8'b00011000;
        13'd2301: m_out<=8'b00010000;
        13'd2302: m_out<=8'b00001110;
        13'd2303: m_out<=8'b00000010;
        13'd2304: m_out<=8'b11111001;
        13'd2305: m_out<=8'b11011111;
        13'd2306: m_out<=8'b11010001;
        13'd2307: m_out<=8'b11111000;
        13'd2308: m_out<=8'b00000100;
        13'd2309: m_out<=8'b11111001;
        13'd2310: m_out<=8'b11101101;
        13'd2311: m_out<=8'b00001101;
        13'd2312: m_out<=8'b00001001;
        13'd2313: m_out<=8'b00111110;
        13'd2314: m_out<=8'b11110111;
        13'd2315: m_out<=8'b00011101;
        13'd2316: m_out<=8'b11010110;
        13'd2317: m_out<=8'b00000010;
        13'd2318: m_out<=8'b00000000;
        13'd2319: m_out<=8'b00100000;
        13'd2320: m_out<=8'b11111010;
        13'd2321: m_out<=8'b00001010;
        13'd2322: m_out<=8'b11111101;
        13'd2323: m_out<=8'b11101100;
        13'd2324: m_out<=8'b11111010;
        13'd2325: m_out<=8'b00011100;
        13'd2326: m_out<=8'b11011001;
        13'd2327: m_out<=8'b00000111;
        13'd2328: m_out<=8'b11111010;
        13'd2329: m_out<=8'b00001000;
        13'd2330: m_out<=8'b00000101;
        13'd2331: m_out<=8'b00000000;
        13'd2332: m_out<=8'b11101000;
        13'd2333: m_out<=8'b11111101;
        13'd2334: m_out<=8'b11101011;
        13'd2335: m_out<=8'b00000011;
        13'd2336: m_out<=8'b11100111;
        13'd2337: m_out<=8'b00010011;
        13'd2338: m_out<=8'b11100001;
        13'd2339: m_out<=8'b00010111;
        13'd2340: m_out<=8'b11100110;
        13'd2341: m_out<=8'b00011110;
        13'd2342: m_out<=8'b11111010;
        13'd2343: m_out<=8'b11101010;
        13'd2344: m_out<=8'b00001110;
        13'd2345: m_out<=8'b11111011;
        13'd2346: m_out<=8'b00000101;
        13'd2347: m_out<=8'b11011011;
        13'd2348: m_out<=8'b11111000;
        13'd2349: m_out<=8'b00011100;
        13'd2350: m_out<=8'b11100110;
        13'd2351: m_out<=8'b10101100;
        13'd2352: m_out<=8'b11011011;
        13'd2353: m_out<=8'b00110010;
        13'd2354: m_out<=8'b11000111;
        13'd2355: m_out<=8'b00010000;
        13'd2356: m_out<=8'b00011011;
        13'd2357: m_out<=8'b00001101;
        13'd2358: m_out<=8'b00100101;
        13'd2359: m_out<=8'b11100010;
        13'd2360: m_out<=8'b00011111;
        13'd2361: m_out<=8'b11111000;
        13'd2362: m_out<=8'b00011110;
        13'd2363: m_out<=8'b11110101;
        13'd2364: m_out<=8'b00100011;
        13'd2365: m_out<=8'b11000100;
        13'd2366: m_out<=8'b00100110;
        13'd2367: m_out<=8'b00001100;
        13'd2368: m_out<=8'b00011111;
        13'd2369: m_out<=8'b11011110;
        13'd2370: m_out<=8'b11111001;
        13'd2371: m_out<=8'b11001001;
        13'd2372: m_out<=8'b11101100;
        13'd2373: m_out<=8'b11010011;
        13'd2374: m_out<=8'b11100111;
        13'd2375: m_out<=8'b11100101;
        13'd2376: m_out<=8'b11101100;
        13'd2377: m_out<=8'b11111000;
        13'd2378: m_out<=8'b11011011;
        13'd2379: m_out<=8'b00000010;
        13'd2380: m_out<=8'b11111110;
        13'd2381: m_out<=8'b11101100;
        13'd2382: m_out<=8'b11111011;
        13'd2383: m_out<=8'b00100110;
        13'd2384: m_out<=8'b11111101;
        13'd2385: m_out<=8'b00001110;
        13'd2386: m_out<=8'b11101101;
        13'd2387: m_out<=8'b00100001;
        13'd2388: m_out<=8'b11110010;
        13'd2389: m_out<=8'b00001000;
        13'd2390: m_out<=8'b11100111;
        13'd2391: m_out<=8'b00000101;
        13'd2392: m_out<=8'b11100100;
        13'd2393: m_out<=8'b00001101;
        13'd2394: m_out<=8'b00000010;
        13'd2395: m_out<=8'b00010000;
        13'd2396: m_out<=8'b00001000;
        13'd2397: m_out<=8'b00100000;
        13'd2398: m_out<=8'b11111101;
        13'd2399: m_out<=8'b11100111;
        13'd2400: m_out<=8'b11011010;
        13'd2401: m_out<=8'b11011101;
        13'd2402: m_out<=8'b11101111;
        13'd2403: m_out<=8'b00000000;
        13'd2404: m_out<=8'b00001000;
        13'd2405: m_out<=8'b11011011;
        13'd2406: m_out<=8'b00100110;
        13'd2407: m_out<=8'b11010000;
        13'd2408: m_out<=8'b00001110;
        13'd2409: m_out<=8'b00001000;
        13'd2410: m_out<=8'b11101110;
        13'd2411: m_out<=8'b11001101;
        13'd2412: m_out<=8'b00001001;
        13'd2413: m_out<=8'b00111001;
        13'd2414: m_out<=8'b00001111;
        13'd2415: m_out<=8'b00010011;
        13'd2416: m_out<=8'b11110000;
        13'd2417: m_out<=8'b11101010;
        13'd2418: m_out<=8'b00000101;
        13'd2419: m_out<=8'b11111001;
        13'd2420: m_out<=8'b00100001;
        13'd2421: m_out<=8'b00011011;
        13'd2422: m_out<=8'b00001011;
        13'd2423: m_out<=8'b00001101;
        13'd2424: m_out<=8'b11110111;
        13'd2425: m_out<=8'b11100110;
        13'd2426: m_out<=8'b00100110;
        13'd2427: m_out<=8'b11100001;
        13'd2428: m_out<=8'b00001010;
        13'd2429: m_out<=8'b11111000;
        13'd2430: m_out<=8'b00000000;
        13'd2431: m_out<=8'b11111010;
        13'd2432: m_out<=8'b11100100;
        13'd2433: m_out<=8'b00010010;
        13'd2434: m_out<=8'b00001001;
        13'd2435: m_out<=8'b00001010;
        13'd2436: m_out<=8'b11011001;
        13'd2437: m_out<=8'b00000111;
        13'd2438: m_out<=8'b11100000;
        13'd2439: m_out<=8'b11101010;
        13'd2440: m_out<=8'b00001111;
        13'd2441: m_out<=8'b00001000;
        13'd2442: m_out<=8'b00011010;
        13'd2443: m_out<=8'b00100110;
        13'd2444: m_out<=8'b11110100;
        13'd2445: m_out<=8'b00001110;
        13'd2446: m_out<=8'b00101110;
        13'd2447: m_out<=8'b11011101;
        13'd2448: m_out<=8'b11100010;
        13'd2449: m_out<=8'b00000110;
        13'd2450: m_out<=8'b00011111;
        13'd2451: m_out<=8'b00011101;
        13'd2452: m_out<=8'b11111110;
        13'd2453: m_out<=8'b00010000;
        13'd2454: m_out<=8'b11101010;
        13'd2455: m_out<=8'b00011010;
        13'd2456: m_out<=8'b00010001;
        13'd2457: m_out<=8'b11110111;
        13'd2458: m_out<=8'b00011100;
        13'd2459: m_out<=8'b00001101;
        13'd2460: m_out<=8'b00101000;
        13'd2461: m_out<=8'b00011011;
        13'd2462: m_out<=8'b11110001;
        13'd2463: m_out<=8'b00101010;
        13'd2464: m_out<=8'b11010101;
        13'd2465: m_out<=8'b11001011;
        13'd2466: m_out<=8'b00010010;
        13'd2467: m_out<=8'b11110100;
        13'd2468: m_out<=8'b11011000;
        13'd2469: m_out<=8'b00010110;
        13'd2470: m_out<=8'b00011111;
        13'd2471: m_out<=8'b11110001;
        13'd2472: m_out<=8'b00000100;
        13'd2473: m_out<=8'b00100011;
        13'd2474: m_out<=8'b00001000;
        13'd2475: m_out<=8'b11001101;
        13'd2476: m_out<=8'b00010111;
        13'd2477: m_out<=8'b00010010;
        13'd2478: m_out<=8'b11010100;
        13'd2479: m_out<=8'b00001001;
        13'd2480: m_out<=8'b00010111;
        13'd2481: m_out<=8'b00001010;
        13'd2482: m_out<=8'b11111101;
        13'd2483: m_out<=8'b00100101;
        13'd2484: m_out<=8'b00101000;
        13'd2485: m_out<=8'b00000110;
        13'd2486: m_out<=8'b00010100;
        13'd2487: m_out<=8'b11111100;
        13'd2488: m_out<=8'b00001001;
        13'd2489: m_out<=8'b11101011;
        13'd2490: m_out<=8'b00001001;
        13'd2491: m_out<=8'b11010011;
        13'd2492: m_out<=8'b11101101;
        13'd2493: m_out<=8'b11111010;
        13'd2494: m_out<=8'b11110111;
        13'd2495: m_out<=8'b00110001;
        13'd2496: m_out<=8'b11011100;
        13'd2497: m_out<=8'b11100011;
        13'd2498: m_out<=8'b11110111;
        13'd2499: m_out<=8'b11110010;
        13'd2500: m_out<=8'b00000000;
        13'd2501: m_out<=8'b11011111;
        13'd2502: m_out<=8'b00010010;
        13'd2503: m_out<=8'b11101000;
        13'd2504: m_out<=8'b11111111;
        13'd2505: m_out<=8'b11101000;
        13'd2506: m_out<=8'b00000000;
        13'd2507: m_out<=8'b00011110;
        13'd2508: m_out<=8'b11101111;
        13'd2509: m_out<=8'b11100101;
        13'd2510: m_out<=8'b11110101;
        13'd2511: m_out<=8'b11111000;
        13'd2512: m_out<=8'b11000010;
        13'd2513: m_out<=8'b00000101;
        13'd2514: m_out<=8'b11101100;
        13'd2515: m_out<=8'b00010100;
        13'd2516: m_out<=8'b00011111;
        13'd2517: m_out<=8'b11111111;
        13'd2518: m_out<=8'b11111100;
        13'd2519: m_out<=8'b11101011;
        13'd2520: m_out<=8'b11111100;
        13'd2521: m_out<=8'b00001001;
        13'd2522: m_out<=8'b11110000;
        13'd2523: m_out<=8'b11111010;
        13'd2524: m_out<=8'b11110101;
        13'd2525: m_out<=8'b11111100;
        13'd2526: m_out<=8'b00000000;
        13'd2527: m_out<=8'b11110000;
        13'd2528: m_out<=8'b11101101;
        13'd2529: m_out<=8'b11111101;
        13'd2530: m_out<=8'b00001111;
        13'd2531: m_out<=8'b11110001;
        13'd2532: m_out<=8'b11111010;
        13'd2533: m_out<=8'b00010000;
        13'd2534: m_out<=8'b11100111;
        13'd2535: m_out<=8'b11110000;
        13'd2536: m_out<=8'b11110011;
        13'd2537: m_out<=8'b11011000;
        13'd2538: m_out<=8'b11111000;
        13'd2539: m_out<=8'b00011110;
        13'd2540: m_out<=8'b11011101;
        13'd2541: m_out<=8'b11101010;
        13'd2542: m_out<=8'b11110011;
        13'd2543: m_out<=8'b11001111;
        13'd2544: m_out<=8'b11110011;
        13'd2545: m_out<=8'b00001111;
        13'd2546: m_out<=8'b00101110;
        13'd2547: m_out<=8'b00011000;
        13'd2548: m_out<=8'b00001010;
        13'd2549: m_out<=8'b00011000;
        13'd2550: m_out<=8'b11101000;
        13'd2551: m_out<=8'b11101100;
        13'd2552: m_out<=8'b11110101;
        13'd2553: m_out<=8'b11100011;
        13'd2554: m_out<=8'b11111101;
        13'd2555: m_out<=8'b11010100;
        13'd2556: m_out<=8'b00000110;
        13'd2557: m_out<=8'b00000011;
        13'd2558: m_out<=8'b00011100;
        13'd2559: m_out<=8'b11110110;
        13'd2560: m_out<=8'b00011011;
        13'd2561: m_out<=8'b00000000;
        13'd2562: m_out<=8'b00001000;
        13'd2563: m_out<=8'b00100101;
        13'd2564: m_out<=8'b01000001;
        13'd2565: m_out<=8'b00101110;
        13'd2566: m_out<=8'b00000000;
        13'd2567: m_out<=8'b00010010;
        13'd2568: m_out<=8'b00000101;
        13'd2569: m_out<=8'b00000001;
        13'd2570: m_out<=8'b11001010;
        13'd2571: m_out<=8'b11111001;
        13'd2572: m_out<=8'b00100111;
        13'd2573: m_out<=8'b00001010;
        13'd2574: m_out<=8'b11101010;
        13'd2575: m_out<=8'b11110101;
        13'd2576: m_out<=8'b00010100;
        13'd2577: m_out<=8'b11101110;
        13'd2578: m_out<=8'b11011011;
        13'd2579: m_out<=8'b11110111;
        13'd2580: m_out<=8'b11100011;
        13'd2581: m_out<=8'b00000000;
        13'd2582: m_out<=8'b01000100;
        13'd2583: m_out<=8'b00010010;
        13'd2584: m_out<=8'b11110100;
        13'd2585: m_out<=8'b00000011;
        13'd2586: m_out<=8'b11100000;
        13'd2587: m_out<=8'b00000011;
        13'd2588: m_out<=8'b00000011;
        13'd2589: m_out<=8'b00100110;
        13'd2590: m_out<=8'b11010111;
        13'd2591: m_out<=8'b11101001;
        13'd2592: m_out<=8'b00001011;
        13'd2593: m_out<=8'b00000111;
        13'd2594: m_out<=8'b00001111;
        13'd2595: m_out<=8'b11010101;
        13'd2596: m_out<=8'b00110100;
        13'd2597: m_out<=8'b00000101;
        13'd2598: m_out<=8'b11101100;
        13'd2599: m_out<=8'b00000010;
        13'd2600: m_out<=8'b00010000;
        13'd2601: m_out<=8'b00001001;
        13'd2602: m_out<=8'b11111101;
        13'd2603: m_out<=8'b11011101;
        13'd2604: m_out<=8'b11100110;
        13'd2605: m_out<=8'b00000101;
        13'd2606: m_out<=8'b00001100;
        13'd2607: m_out<=8'b00001010;
        13'd2608: m_out<=8'b00010110;
        13'd2609: m_out<=8'b00000110;
        13'd2610: m_out<=8'b00001001;
        13'd2611: m_out<=8'b11101011;
        13'd2612: m_out<=8'b00000011;
        13'd2613: m_out<=8'b00000011;
        13'd2614: m_out<=8'b00100100;
        13'd2615: m_out<=8'b00100001;
        13'd2616: m_out<=8'b00011101;
        13'd2617: m_out<=8'b00001011;
        13'd2618: m_out<=8'b11111001;
        13'd2619: m_out<=8'b11111001;
        13'd2620: m_out<=8'b00000010;
        13'd2621: m_out<=8'b00010001;
        13'd2622: m_out<=8'b11111110;
        13'd2623: m_out<=8'b11110001;
        13'd2624: m_out<=8'b00011101;
        13'd2625: m_out<=8'b11111011;
        13'd2626: m_out<=8'b11110110;
        13'd2627: m_out<=8'b11100011;
        13'd2628: m_out<=8'b11111000;
        13'd2629: m_out<=8'b11110011;
        13'd2630: m_out<=8'b11100100;
        13'd2631: m_out<=8'b00010101;
        13'd2632: m_out<=8'b00011101;
        13'd2633: m_out<=8'b11010100;
        13'd2634: m_out<=8'b11110101;
        13'd2635: m_out<=8'b00001001;
        13'd2636: m_out<=8'b00000011;
        13'd2637: m_out<=8'b11001111;
        13'd2638: m_out<=8'b11100001;
        13'd2639: m_out<=8'b00010010;
        13'd2640: m_out<=8'b00000001;
        13'd2641: m_out<=8'b11111010;
        13'd2642: m_out<=8'b00000011;
        13'd2643: m_out<=8'b00010011;
        13'd2644: m_out<=8'b00001001;
        13'd2645: m_out<=8'b00010000;
        13'd2646: m_out<=8'b00001000;
        13'd2647: m_out<=8'b11111110;
        13'd2648: m_out<=8'b00010100;
        13'd2649: m_out<=8'b00001100;
        13'd2650: m_out<=8'b00011010;
        13'd2651: m_out<=8'b00000101;
        13'd2652: m_out<=8'b11110111;
        13'd2653: m_out<=8'b11010011;
        13'd2654: m_out<=8'b11110100;
        13'd2655: m_out<=8'b11101101;
        13'd2656: m_out<=8'b11101001;
        13'd2657: m_out<=8'b00000010;
        13'd2658: m_out<=8'b11110110;
        13'd2659: m_out<=8'b00010011;
        13'd2660: m_out<=8'b11011110;
        13'd2661: m_out<=8'b11110111;
        13'd2662: m_out<=8'b11110111;
        13'd2663: m_out<=8'b11011100;
        13'd2664: m_out<=8'b10111111;
        13'd2665: m_out<=8'b00001001;
        13'd2666: m_out<=8'b00110110;
        13'd2667: m_out<=8'b01000100;
        13'd2668: m_out<=8'b11111111;
        13'd2669: m_out<=8'b11001000;
        13'd2670: m_out<=8'b11110000;
        13'd2671: m_out<=8'b00001100;
        13'd2672: m_out<=8'b00001111;
        13'd2673: m_out<=8'b00001110;
        13'd2674: m_out<=8'b11110011;
        13'd2675: m_out<=8'b00011001;
        13'd2676: m_out<=8'b11011011;
        13'd2677: m_out<=8'b00000010;
        13'd2678: m_out<=8'b11100010;
        13'd2679: m_out<=8'b11101110;
        13'd2680: m_out<=8'b11111111;
        13'd2681: m_out<=8'b00010100;
        13'd2682: m_out<=8'b00000000;
        13'd2683: m_out<=8'b11101100;
        13'd2684: m_out<=8'b11101001;
        13'd2685: m_out<=8'b00110011;
        13'd2686: m_out<=8'b00100110;
        13'd2687: m_out<=8'b00110111;
        13'd2688: m_out<=8'b11011001;
        13'd2689: m_out<=8'b11111001;
        13'd2690: m_out<=8'b11100011;
        13'd2691: m_out<=8'b00000100;
        13'd2692: m_out<=8'b00011100;
        13'd2693: m_out<=8'b00011000;
        13'd2694: m_out<=8'b01000100;
        13'd2695: m_out<=8'b11110011;
        13'd2696: m_out<=8'b00000011;
        13'd2697: m_out<=8'b00011111;
        13'd2698: m_out<=8'b00010111;
        13'd2699: m_out<=8'b00000001;
        13'd2700: m_out<=8'b11110001;
        13'd2701: m_out<=8'b11111101;
        13'd2702: m_out<=8'b11111011;
        13'd2703: m_out<=8'b00000101;
        13'd2704: m_out<=8'b11100110;
        13'd2705: m_out<=8'b00100101;
        13'd2706: m_out<=8'b00000111;
        13'd2707: m_out<=8'b11110000;
        13'd2708: m_out<=8'b00010000;
        13'd2709: m_out<=8'b00001110;
        13'd2710: m_out<=8'b00011011;
        13'd2711: m_out<=8'b00000010;
        13'd2712: m_out<=8'b00001101;
        13'd2713: m_out<=8'b11100001;
        13'd2714: m_out<=8'b11110001;
        13'd2715: m_out<=8'b11111010;
        13'd2716: m_out<=8'b00001100;
        13'd2717: m_out<=8'b00101011;
        13'd2718: m_out<=8'b11101000;
        13'd2719: m_out<=8'b00001110;
        13'd2720: m_out<=8'b00010110;
        13'd2721: m_out<=8'b00000100;
        13'd2722: m_out<=8'b11111010;
        13'd2723: m_out<=8'b11111001;
        13'd2724: m_out<=8'b00110010;
        13'd2725: m_out<=8'b00000001;
        13'd2726: m_out<=8'b00100111;
        13'd2727: m_out<=8'b00011111;
        13'd2728: m_out<=8'b00100010;
        13'd2729: m_out<=8'b00010111;
        13'd2730: m_out<=8'b00010010;
        13'd2731: m_out<=8'b11110001;
        13'd2732: m_out<=8'b00100110;
        13'd2733: m_out<=8'b00000011;
        13'd2734: m_out<=8'b00001110;
        13'd2735: m_out<=8'b11011101;
        13'd2736: m_out<=8'b00010010;
        13'd2737: m_out<=8'b11110110;
        13'd2738: m_out<=8'b11011001;
        13'd2739: m_out<=8'b11101100;
        13'd2740: m_out<=8'b11110111;
        13'd2741: m_out<=8'b00000001;
        13'd2742: m_out<=8'b00101101;
        13'd2743: m_out<=8'b00111000;
        13'd2744: m_out<=8'b00111011;
        13'd2745: m_out<=8'b00011110;
        13'd2746: m_out<=8'b11011100;
        13'd2747: m_out<=8'b00000100;
        13'd2748: m_out<=8'b00010101;
        13'd2749: m_out<=8'b00010001;
        13'd2750: m_out<=8'b00011010;
        13'd2751: m_out<=8'b00011101;
        13'd2752: m_out<=8'b11101100;
        13'd2753: m_out<=8'b11101000;
        13'd2754: m_out<=8'b00000101;
        13'd2755: m_out<=8'b00011010;
        13'd2756: m_out<=8'b00001110;
        13'd2757: m_out<=8'b00110111;
        13'd2758: m_out<=8'b11011111;
        13'd2759: m_out<=8'b00001001;
        13'd2760: m_out<=8'b11000101;
        13'd2761: m_out<=8'b11111011;
        13'd2762: m_out<=8'b00100110;
        13'd2763: m_out<=8'b11111100;
        13'd2764: m_out<=8'b00010100;
        13'd2765: m_out<=8'b11010001;
        13'd2766: m_out<=8'b11101010;
        13'd2767: m_out<=8'b11110000;
        13'd2768: m_out<=8'b11101111;
        13'd2769: m_out<=8'b00001011;
        13'd2770: m_out<=8'b00001010;
        13'd2771: m_out<=8'b00110101;
        13'd2772: m_out<=8'b01000000;
        13'd2773: m_out<=8'b00100010;
        13'd2774: m_out<=8'b11111110;
        13'd2775: m_out<=8'b00101010;
        13'd2776: m_out<=8'b11101110;
        13'd2777: m_out<=8'b00010101;
        13'd2778: m_out<=8'b11100100;
        13'd2779: m_out<=8'b11110001;
        13'd2780: m_out<=8'b11100100;
        13'd2781: m_out<=8'b00101111;
        13'd2782: m_out<=8'b11101000;
        13'd2783: m_out<=8'b11100111;
        13'd2784: m_out<=8'b00001110;
        13'd2785: m_out<=8'b00110100;
        13'd2786: m_out<=8'b11110000;
        13'd2787: m_out<=8'b00100111;
        13'd2788: m_out<=8'b00011001;
        13'd2789: m_out<=8'b00010011;
        13'd2790: m_out<=8'b11001111;
        13'd2791: m_out<=8'b11110100;
        13'd2792: m_out<=8'b11111000;
        13'd2793: m_out<=8'b11111111;
        13'd2794: m_out<=8'b11111000;
        13'd2795: m_out<=8'b11111001;
        13'd2796: m_out<=8'b11111001;
        13'd2797: m_out<=8'b11110110;
        13'd2798: m_out<=8'b00101010;
        13'd2799: m_out<=8'b00001100;
        13'd2800: m_out<=8'b00011011;
        13'd2801: m_out<=8'b00001011;
        13'd2802: m_out<=8'b11101010;
        13'd2803: m_out<=8'b11111000;
        13'd2804: m_out<=8'b00010110;
        13'd2805: m_out<=8'b00000101;
        13'd2806: m_out<=8'b00000000;
        13'd2807: m_out<=8'b11111000;
        13'd2808: m_out<=8'b00010100;
        13'd2809: m_out<=8'b00010001;
        13'd2810: m_out<=8'b11011010;
        13'd2811: m_out<=8'b00011101;
        13'd2812: m_out<=8'b00111110;
        13'd2813: m_out<=8'b00000010;
        13'd2814: m_out<=8'b11101110;
        13'd2815: m_out<=8'b00000111;
        13'd2816: m_out<=8'b11100100;
        13'd2817: m_out<=8'b00001010;
        13'd2818: m_out<=8'b00001010;
        13'd2819: m_out<=8'b11110110;
        13'd2820: m_out<=8'b11011011;
        13'd2821: m_out<=8'b00110100;
        13'd2822: m_out<=8'b00011000;
        13'd2823: m_out<=8'b00100100;
        13'd2824: m_out<=8'b11111100;
        13'd2825: m_out<=8'b11111011;
        13'd2826: m_out<=8'b00000011;
        13'd2827: m_out<=8'b00101010;
        13'd2828: m_out<=8'b11011110;
        13'd2829: m_out<=8'b11101100;
        13'd2830: m_out<=8'b00000110;
        13'd2831: m_out<=8'b11101100;
        13'd2832: m_out<=8'b00011001;
        13'd2833: m_out<=8'b11111000;
        13'd2834: m_out<=8'b00001001;
        13'd2835: m_out<=8'b00001010;
        13'd2836: m_out<=8'b00000101;
        13'd2837: m_out<=8'b00000001;
        13'd2838: m_out<=8'b11110001;
        13'd2839: m_out<=8'b00010000;
        13'd2840: m_out<=8'b00001111;
        13'd2841: m_out<=8'b11011111;
        13'd2842: m_out<=8'b11110001;
        13'd2843: m_out<=8'b11000011;
        13'd2844: m_out<=8'b00001100;
        13'd2845: m_out<=8'b11110100;
        13'd2846: m_out<=8'b11111010;
        13'd2847: m_out<=8'b00100011;
        13'd2848: m_out<=8'b00011100;
        13'd2849: m_out<=8'b11011101;
        13'd2850: m_out<=8'b00000001;
        13'd2851: m_out<=8'b00001001;
        13'd2852: m_out<=8'b11100101;
        13'd2853: m_out<=8'b11101010;
        13'd2854: m_out<=8'b00011100;
        13'd2855: m_out<=8'b11101010;
        13'd2856: m_out<=8'b11111101;
        13'd2857: m_out<=8'b00110010;
        13'd2858: m_out<=8'b11110111;
        13'd2859: m_out<=8'b11110000;
        13'd2860: m_out<=8'b11010101;
        13'd2861: m_out<=8'b00000001;
        13'd2862: m_out<=8'b00010100;
        13'd2863: m_out<=8'b00011010;
        13'd2864: m_out<=8'b11101010;
        13'd2865: m_out<=8'b00000011;
        13'd2866: m_out<=8'b00011000;
        13'd2867: m_out<=8'b00011000;
        13'd2868: m_out<=8'b11110011;
        13'd2869: m_out<=8'b00100001;
        13'd2870: m_out<=8'b00011101;
        13'd2871: m_out<=8'b00111001;
        13'd2872: m_out<=8'b00001000;
        13'd2873: m_out<=8'b11110000;
        13'd2874: m_out<=8'b00100000;
        13'd2875: m_out<=8'b00001001;
        13'd2876: m_out<=8'b11100000;
        13'd2877: m_out<=8'b00100000;
        13'd2878: m_out<=8'b00000011;
        13'd2879: m_out<=8'b00001111;
        13'd2880: m_out<=8'b11101110;
        13'd2881: m_out<=8'b00000001;
        13'd2882: m_out<=8'b00000010;
        13'd2883: m_out<=8'b00001111;
        13'd2884: m_out<=8'b11011011;
        13'd2885: m_out<=8'b00000101;
        13'd2886: m_out<=8'b11111011;
        13'd2887: m_out<=8'b00000000;
        13'd2888: m_out<=8'b11101011;
        13'd2889: m_out<=8'b11011111;
        13'd2890: m_out<=8'b00010001;
        13'd2891: m_out<=8'b00010110;
        13'd2892: m_out<=8'b11110110;
        13'd2893: m_out<=8'b11110001;
        13'd2894: m_out<=8'b00001001;
        13'd2895: m_out<=8'b00001010;
        13'd2896: m_out<=8'b11101001;
        13'd2897: m_out<=8'b00011000;
        13'd2898: m_out<=8'b00010011;
        13'd2899: m_out<=8'b11010100;
        13'd2900: m_out<=8'b00000010;
        13'd2901: m_out<=8'b00100000;
        13'd2902: m_out<=8'b00000110;
        13'd2903: m_out<=8'b00011100;
        13'd2904: m_out<=8'b11110111;
        13'd2905: m_out<=8'b00100001;
        13'd2906: m_out<=8'b11100101;
        13'd2907: m_out<=8'b00011000;
        13'd2908: m_out<=8'b00000101;
        13'd2909: m_out<=8'b11101011;
        13'd2910: m_out<=8'b00010001;
        13'd2911: m_out<=8'b00011011;
        13'd2912: m_out<=8'b11100010;
        13'd2913: m_out<=8'b00000010;
        13'd2914: m_out<=8'b11101010;
        13'd2915: m_out<=8'b00001011;
        13'd2916: m_out<=8'b11101111;
        13'd2917: m_out<=8'b11001101;
        13'd2918: m_out<=8'b00001100;
        13'd2919: m_out<=8'b10111100;
        13'd2920: m_out<=8'b11110110;
        13'd2921: m_out<=8'b11101001;
        13'd2922: m_out<=8'b00011100;
        13'd2923: m_out<=8'b00010001;
        13'd2924: m_out<=8'b00110011;
        13'd2925: m_out<=8'b00000101;
        13'd2926: m_out<=8'b00010110;
        13'd2927: m_out<=8'b00011110;
        13'd2928: m_out<=8'b11110011;
        13'd2929: m_out<=8'b11111010;
        13'd2930: m_out<=8'b11101111;
        13'd2931: m_out<=8'b11001001;
        13'd2932: m_out<=8'b00000111;
        13'd2933: m_out<=8'b00010101;
        13'd2934: m_out<=8'b00001011;
        13'd2935: m_out<=8'b00001001;
        13'd2936: m_out<=8'b11110101;
        13'd2937: m_out<=8'b11000000;
        13'd2938: m_out<=8'b00010110;
        13'd2939: m_out<=8'b00001100;
        13'd2940: m_out<=8'b00000100;
        13'd2941: m_out<=8'b11100101;
        13'd2942: m_out<=8'b11110011;
        13'd2943: m_out<=8'b00010110;
        13'd2944: m_out<=8'b00001010;
        13'd2945: m_out<=8'b11001011;
        13'd2946: m_out<=8'b11001011;
        13'd2947: m_out<=8'b11111111;
        13'd2948: m_out<=8'b00100101;
        13'd2949: m_out<=8'b11101001;
        13'd2950: m_out<=8'b00110100;
        13'd2951: m_out<=8'b11111000;
        13'd2952: m_out<=8'b11100110;
        13'd2953: m_out<=8'b11101001;
        13'd2954: m_out<=8'b00001000;
        13'd2955: m_out<=8'b00011001;
        13'd2956: m_out<=8'b11100110;
        13'd2957: m_out<=8'b00100101;
        13'd2958: m_out<=8'b00010100;
        13'd2959: m_out<=8'b11101010;
        13'd2960: m_out<=8'b11101111;
        13'd2961: m_out<=8'b10111101;
        13'd2962: m_out<=8'b00010100;
        13'd2963: m_out<=8'b00000011;
        13'd2964: m_out<=8'b00011011;
        13'd2965: m_out<=8'b11100100;
        13'd2966: m_out<=8'b11101110;
        13'd2967: m_out<=8'b11101101;
        13'd2968: m_out<=8'b11110101;
        13'd2969: m_out<=8'b11011111;
        13'd2970: m_out<=8'b00010011;
        13'd2971: m_out<=8'b00110011;
        13'd2972: m_out<=8'b11101101;
        13'd2973: m_out<=8'b00001001;
        13'd2974: m_out<=8'b00000010;
        13'd2975: m_out<=8'b11101100;
        13'd2976: m_out<=8'b00100000;
        13'd2977: m_out<=8'b00100001;
        13'd2978: m_out<=8'b00001000;
        13'd2979: m_out<=8'b00011011;
        13'd2980: m_out<=8'b00010101;
        13'd2981: m_out<=8'b11100111;
        13'd2982: m_out<=8'b00011010;
        13'd2983: m_out<=8'b00000000;
        13'd2984: m_out<=8'b00010011;
        13'd2985: m_out<=8'b00010111;
        13'd2986: m_out<=8'b11111001;
        13'd2987: m_out<=8'b11101111;
        13'd2988: m_out<=8'b00000111;
        13'd2989: m_out<=8'b00010101;
        13'd2990: m_out<=8'b00000101;
        13'd2991: m_out<=8'b11111001;
        13'd2992: m_out<=8'b00000001;
        13'd2993: m_out<=8'b11110011;
        13'd2994: m_out<=8'b00111010;
        13'd2995: m_out<=8'b11011111;
        13'd2996: m_out<=8'b11100000;
        13'd2997: m_out<=8'b11110111;
        13'd2998: m_out<=8'b11110010;
        13'd2999: m_out<=8'b00001101;
        13'd3000: m_out<=8'b00011101;
        13'd3001: m_out<=8'b00001100;
        13'd3002: m_out<=8'b00000101;
        13'd3003: m_out<=8'b00101011;
        13'd3004: m_out<=8'b01000111;
        13'd3005: m_out<=8'b01010100;
        13'd3006: m_out<=8'b00000011;
        13'd3007: m_out<=8'b01000011;
        13'd3008: m_out<=8'b00010110;
        13'd3009: m_out<=8'b00001011;
        13'd3010: m_out<=8'b00101001;
        13'd3011: m_out<=8'b11001111;
        13'd3012: m_out<=8'b00001010;
        13'd3013: m_out<=8'b11010000;
        13'd3014: m_out<=8'b10011111;
        13'd3015: m_out<=8'b10011111;
        13'd3016: m_out<=8'b11011110;
        13'd3017: m_out<=8'b10111101;
        13'd3018: m_out<=8'b10100010;
        13'd3019: m_out<=8'b11010100;
        13'd3020: m_out<=8'b11111001;
        13'd3021: m_out<=8'b11111101;
        13'd3022: m_out<=8'b11111101;
        13'd3023: m_out<=8'b00001011;
        13'd3024: m_out<=8'b11110010;
        13'd3025: m_out<=8'b00000001;
        13'd3026: m_out<=8'b11111010;
        13'd3027: m_out<=8'b00010000;
        13'd3028: m_out<=8'b00001101;
        13'd3029: m_out<=8'b11110100;
        13'd3030: m_out<=8'b00101111;
        13'd3031: m_out<=8'b11100000;
        13'd3032: m_out<=8'b00111010;
        13'd3033: m_out<=8'b00011001;
        13'd3034: m_out<=8'b00010000;
        13'd3035: m_out<=8'b11111110;
        13'd3036: m_out<=8'b00010110;
        13'd3037: m_out<=8'b00011011;
        13'd3038: m_out<=8'b11100100;
        13'd3039: m_out<=8'b11101100;
        13'd3040: m_out<=8'b11111100;
        13'd3041: m_out<=8'b00010100;
        13'd3042: m_out<=8'b00100000;
        13'd3043: m_out<=8'b00000001;
        13'd3044: m_out<=8'b11101010;
        13'd3045: m_out<=8'b11101001;
        13'd3046: m_out<=8'b00001011;
        13'd3047: m_out<=8'b11100111;
        13'd3048: m_out<=8'b00011100;
        13'd3049: m_out<=8'b00000000;
        13'd3050: m_out<=8'b11110111;
        13'd3051: m_out<=8'b00100100;
        13'd3052: m_out<=8'b11100110;
        13'd3053: m_out<=8'b00011010;
        13'd3054: m_out<=8'b11101001;
        13'd3055: m_out<=8'b11101000;
        13'd3056: m_out<=8'b00000101;
        13'd3057: m_out<=8'b00000100;
        13'd3058: m_out<=8'b11101011;
        13'd3059: m_out<=8'b11110100;
        13'd3060: m_out<=8'b11100000;
        13'd3061: m_out<=8'b11100011;
        13'd3062: m_out<=8'b00000101;
        13'd3063: m_out<=8'b11101001;
        13'd3064: m_out<=8'b11011111;
        13'd3065: m_out<=8'b11011001;
        13'd3066: m_out<=8'b11110111;
        13'd3067: m_out<=8'b11111001;
        13'd3068: m_out<=8'b11100010;
        13'd3069: m_out<=8'b11011011;
        13'd3070: m_out<=8'b00000101;
        13'd3071: m_out<=8'b00001111;
        13'd3072: m_out<=8'b11110100;
        13'd3073: m_out<=8'b11111111;
        13'd3074: m_out<=8'b00011011;
        13'd3075: m_out<=8'b11100010;
        13'd3076: m_out<=8'b11111011;
        13'd3077: m_out<=8'b00001010;
        13'd3078: m_out<=8'b00001011;
        13'd3079: m_out<=8'b00010011;
        13'd3080: m_out<=8'b11101101;
        13'd3081: m_out<=8'b11101010;
        13'd3082: m_out<=8'b11111010;
        13'd3083: m_out<=8'b00000001;
        13'd3084: m_out<=8'b11100111;
        13'd3085: m_out<=8'b00101001;
        13'd3086: m_out<=8'b10111100;
        13'd3087: m_out<=8'b00011001;
        13'd3088: m_out<=8'b00011111;
        13'd3089: m_out<=8'b00100011;
        13'd3090: m_out<=8'b11111011;
        13'd3091: m_out<=8'b00001001;
        13'd3092: m_out<=8'b11100110;
        13'd3093: m_out<=8'b00100001;
        13'd3094: m_out<=8'b00100011;
        13'd3095: m_out<=8'b00011101;
        13'd3096: m_out<=8'b00000111;
        13'd3097: m_out<=8'b11100111;
        13'd3098: m_out<=8'b00100110;
        13'd3099: m_out<=8'b00001111;
        13'd3100: m_out<=8'b00000110;
        13'd3101: m_out<=8'b11011101;
        13'd3102: m_out<=8'b00001100;
        13'd3103: m_out<=8'b11111101;
        13'd3104: m_out<=8'b11111101;
        13'd3105: m_out<=8'b00001011;
        13'd3106: m_out<=8'b11101111;
        13'd3107: m_out<=8'b11111010;
        13'd3108: m_out<=8'b11010110;
        13'd3109: m_out<=8'b00101001;
        13'd3110: m_out<=8'b00101010;
        13'd3111: m_out<=8'b00011100;
        13'd3112: m_out<=8'b00010001;
        13'd3113: m_out<=8'b11011111;
        13'd3114: m_out<=8'b11110110;
        13'd3115: m_out<=8'b00010010;
        13'd3116: m_out<=8'b11100101;
        13'd3117: m_out<=8'b11100011;
        13'd3118: m_out<=8'b11001111;
        13'd3119: m_out<=8'b00001001;
        13'd3120: m_out<=8'b00100010;
        13'd3121: m_out<=8'b11111110;
        13'd3122: m_out<=8'b00000110;
        13'd3123: m_out<=8'b00001000;
        13'd3124: m_out<=8'b11110010;
        13'd3125: m_out<=8'b00000010;
        13'd3126: m_out<=8'b11110001;
        13'd3127: m_out<=8'b11111000;
        13'd3128: m_out<=8'b00001001;
        13'd3129: m_out<=8'b11101111;
        13'd3130: m_out<=8'b00101101;
        13'd3131: m_out<=8'b00001001;
        13'd3132: m_out<=8'b00000111;
        13'd3133: m_out<=8'b11101110;
        13'd3134: m_out<=8'b11110100;
        13'd3135: m_out<=8'b11101001;
        13'd3136: m_out<=8'b00001011;
        13'd3137: m_out<=8'b11110011;
        13'd3138: m_out<=8'b00011000;
        13'd3139: m_out<=8'b00010010;
        13'd3140: m_out<=8'b11111010;
        13'd3141: m_out<=8'b00000000;
        13'd3142: m_out<=8'b00011001;
        13'd3143: m_out<=8'b00110010;
        13'd3144: m_out<=8'b00000001;
        13'd3145: m_out<=8'b11100001;
        13'd3146: m_out<=8'b00001000;
        13'd3147: m_out<=8'b00001000;
        13'd3148: m_out<=8'b11110100;
        13'd3149: m_out<=8'b11011111;
        13'd3150: m_out<=8'b00010101;
        13'd3151: m_out<=8'b00001010;
        13'd3152: m_out<=8'b11101100;
        13'd3153: m_out<=8'b11101000;
        13'd3154: m_out<=8'b11101110;
        13'd3155: m_out<=8'b11000011;
        13'd3156: m_out<=8'b00000010;
        13'd3157: m_out<=8'b00010110;
        13'd3158: m_out<=8'b11111110;
        13'd3159: m_out<=8'b00001100;
        13'd3160: m_out<=8'b00000110;
        13'd3161: m_out<=8'b00011110;
        13'd3162: m_out<=8'b11111111;
        13'd3163: m_out<=8'b00000111;
        13'd3164: m_out<=8'b00010000;
        13'd3165: m_out<=8'b00011001;
        13'd3166: m_out<=8'b00001100;
        13'd3167: m_out<=8'b00011011;
        13'd3168: m_out<=8'b00001101;
        13'd3169: m_out<=8'b00011001;
        13'd3170: m_out<=8'b11111010;
        13'd3171: m_out<=8'b11100100;
        13'd3172: m_out<=8'b11101001;
        13'd3173: m_out<=8'b11100111;
        13'd3174: m_out<=8'b11101110;
        13'd3175: m_out<=8'b00001001;
        13'd3176: m_out<=8'b00110100;
        13'd3177: m_out<=8'b00000010;
        13'd3178: m_out<=8'b00011110;
        13'd3179: m_out<=8'b00000111;
        13'd3180: m_out<=8'b11010011;
        13'd3181: m_out<=8'b11101101;
        13'd3182: m_out<=8'b11110001;
        13'd3183: m_out<=8'b11111111;
        13'd3184: m_out<=8'b00001110;
        13'd3185: m_out<=8'b11011011;
        13'd3186: m_out<=8'b11000111;
        13'd3187: m_out<=8'b00110011;
        13'd3188: m_out<=8'b00001110;
        13'd3189: m_out<=8'b00011101;
        13'd3190: m_out<=8'b00100111;
        13'd3191: m_out<=8'b00001110;
        13'd3192: m_out<=8'b00100001;
        13'd3193: m_out<=8'b11011111;
        13'd3194: m_out<=8'b11111010;
        13'd3195: m_out<=8'b00001100;
        13'd3196: m_out<=8'b11100111;
        13'd3197: m_out<=8'b00001111;
        13'd3198: m_out<=8'b00010101;
        13'd3199: m_out<=8'b11110001;
        13'd3200: m_out<=8'b00010000;
        13'd3201: m_out<=8'b00001000;
        13'd3202: m_out<=8'b11101001;
        13'd3203: m_out<=8'b11110011;
        13'd3204: m_out<=8'b11100111;
        13'd3205: m_out<=8'b00010011;
        13'd3206: m_out<=8'b00011111;
        13'd3207: m_out<=8'b11110111;
        13'd3208: m_out<=8'b11111110;
        13'd3209: m_out<=8'b00000011;
        13'd3210: m_out<=8'b11111111;
        13'd3211: m_out<=8'b00100001;
        13'd3212: m_out<=8'b00110101;
        13'd3213: m_out<=8'b00001010;
        13'd3214: m_out<=8'b11101111;
        13'd3215: m_out<=8'b00001010;
        13'd3216: m_out<=8'b11111100;
        13'd3217: m_out<=8'b00000100;
        13'd3218: m_out<=8'b11111110;
        13'd3219: m_out<=8'b11110010;
        13'd3220: m_out<=8'b11110100;
        13'd3221: m_out<=8'b00000110;
        13'd3222: m_out<=8'b00100111;
        13'd3223: m_out<=8'b00000010;
        13'd3224: m_out<=8'b00000101;
        13'd3225: m_out<=8'b00000001;
        13'd3226: m_out<=8'b11110111;
        13'd3227: m_out<=8'b11101101;
        13'd3228: m_out<=8'b11101100;
        13'd3229: m_out<=8'b11110100;
        13'd3230: m_out<=8'b11010100;
        13'd3231: m_out<=8'b00000101;
        13'd3232: m_out<=8'b11110110;
        13'd3233: m_out<=8'b11100111;
        13'd3234: m_out<=8'b11111000;
        13'd3235: m_out<=8'b00010001;
        13'd3236: m_out<=8'b00010000;
        13'd3237: m_out<=8'b11111010;
        13'd3238: m_out<=8'b11100001;
        13'd3239: m_out<=8'b11101001;
        13'd3240: m_out<=8'b11101110;
        13'd3241: m_out<=8'b00000001;
        13'd3242: m_out<=8'b11111010;
        13'd3243: m_out<=8'b00000100;
        13'd3244: m_out<=8'b11001010;
        13'd3245: m_out<=8'b00000011;
        13'd3246: m_out<=8'b11111111;
        13'd3247: m_out<=8'b00011000;
        13'd3248: m_out<=8'b11111001;
        13'd3249: m_out<=8'b00011000;
        13'd3250: m_out<=8'b11011011;
        13'd3251: m_out<=8'b11001111;
        13'd3252: m_out<=8'b00000101;
        13'd3253: m_out<=8'b11100010;
        13'd3254: m_out<=8'b11110011;
        13'd3255: m_out<=8'b00100101;
        13'd3256: m_out<=8'b00010101;
        13'd3257: m_out<=8'b11011110;
        13'd3258: m_out<=8'b00101110;
        13'd3259: m_out<=8'b00110100;
        13'd3260: m_out<=8'b00000101;
        13'd3261: m_out<=8'b11100010;
        13'd3262: m_out<=8'b00010000;
        13'd3263: m_out<=8'b00001011;
        13'd3264: m_out<=8'b11011110;
        13'd3265: m_out<=8'b00110101;
        13'd3266: m_out<=8'b00000010;
        13'd3267: m_out<=8'b11011001;
        13'd3268: m_out<=8'b00010001;
        13'd3269: m_out<=8'b00010101;
        13'd3270: m_out<=8'b00001101;
        13'd3271: m_out<=8'b00101101;
        13'd3272: m_out<=8'b11100001;
        13'd3273: m_out<=8'b00100000;
        13'd3274: m_out<=8'b00010100;
        13'd3275: m_out<=8'b00001010;
        13'd3276: m_out<=8'b11101010;
        13'd3277: m_out<=8'b11111101;
        13'd3278: m_out<=8'b00001101;
        13'd3279: m_out<=8'b00011100;
        13'd3280: m_out<=8'b11100110;
        13'd3281: m_out<=8'b11101001;
        13'd3282: m_out<=8'b11111101;
        13'd3283: m_out<=8'b00010010;
        13'd3284: m_out<=8'b11100100;
        13'd3285: m_out<=8'b11110111;
        13'd3286: m_out<=8'b01000000;
        13'd3287: m_out<=8'b00001100;
        13'd3288: m_out<=8'b11110101;
        13'd3289: m_out<=8'b11110110;
        13'd3290: m_out<=8'b00101101;
        13'd3291: m_out<=8'b00100010;
        13'd3292: m_out<=8'b11101000;
        13'd3293: m_out<=8'b00011101;
        13'd3294: m_out<=8'b00001100;
        13'd3295: m_out<=8'b11110100;
        13'd3296: m_out<=8'b11111000;
        13'd3297: m_out<=8'b11100000;
        13'd3298: m_out<=8'b11111010;
        13'd3299: m_out<=8'b11100110;
        13'd3300: m_out<=8'b00001001;
        13'd3301: m_out<=8'b11110011;
        13'd3302: m_out<=8'b00001001;
        13'd3303: m_out<=8'b00000001;
        13'd3304: m_out<=8'b11011001;
        13'd3305: m_out<=8'b00011001;
        13'd3306: m_out<=8'b00101100;
        13'd3307: m_out<=8'b00110001;
        13'd3308: m_out<=8'b11110100;
        13'd3309: m_out<=8'b00001010;
        13'd3310: m_out<=8'b11111000;
        13'd3311: m_out<=8'b00000010;
        13'd3312: m_out<=8'b00100000;
        13'd3313: m_out<=8'b00101011;
        13'd3314: m_out<=8'b11101011;
        13'd3315: m_out<=8'b11110101;
        13'd3316: m_out<=8'b11001011;
        13'd3317: m_out<=8'b00001101;
        13'd3318: m_out<=8'b11111101;
        13'd3319: m_out<=8'b11011101;
        13'd3320: m_out<=8'b00000000;
        13'd3321: m_out<=8'b00000010;
        13'd3322: m_out<=8'b11101001;
        13'd3323: m_out<=8'b01000110;
        13'd3324: m_out<=8'b11111010;
        13'd3325: m_out<=8'b00010010;
        13'd3326: m_out<=8'b00001010;
        13'd3327: m_out<=8'b11111100;
        13'd3328: m_out<=8'b00001100;
        13'd3329: m_out<=8'b11110101;
        13'd3330: m_out<=8'b11101010;
        13'd3331: m_out<=8'b01000011;
        13'd3332: m_out<=8'b00000101;
        13'd3333: m_out<=8'b11110001;
        13'd3334: m_out<=8'b00010010;
        13'd3335: m_out<=8'b11010111;
        13'd3336: m_out<=8'b11101111;
        13'd3337: m_out<=8'b11100101;
        13'd3338: m_out<=8'b11110001;
        13'd3339: m_out<=8'b11111101;
        13'd3340: m_out<=8'b11111000;
        13'd3341: m_out<=8'b00111101;
        13'd3342: m_out<=8'b11110110;
        13'd3343: m_out<=8'b11010111;
        13'd3344: m_out<=8'b11010101;
        13'd3345: m_out<=8'b11011111;
        13'd3346: m_out<=8'b00011010;
        13'd3347: m_out<=8'b00100111;
        13'd3348: m_out<=8'b00000101;
        13'd3349: m_out<=8'b00000101;
        13'd3350: m_out<=8'b00100110;
        13'd3351: m_out<=8'b11011010;
        13'd3352: m_out<=8'b00000010;
        13'd3353: m_out<=8'b00010101;
        13'd3354: m_out<=8'b00010001;
        13'd3355: m_out<=8'b11010010;
        13'd3356: m_out<=8'b11111100;
        13'd3357: m_out<=8'b00001111;
        13'd3358: m_out<=8'b00011110;
        13'd3359: m_out<=8'b00000101;
        13'd3360: m_out<=8'b00010001;
        13'd3361: m_out<=8'b00010010;
        13'd3362: m_out<=8'b11011001;
        13'd3363: m_out<=8'b00001101;
        13'd3364: m_out<=8'b11100101;
        13'd3365: m_out<=8'b11110110;
        13'd3366: m_out<=8'b00011001;
        13'd3367: m_out<=8'b11101010;
        13'd3368: m_out<=8'b11111011;
        13'd3369: m_out<=8'b11100001;
        13'd3370: m_out<=8'b00110101;
        13'd3371: m_out<=8'b11101000;
        13'd3372: m_out<=8'b00010011;
        13'd3373: m_out<=8'b01000101;
        13'd3374: m_out<=8'b11101011;
        13'd3375: m_out<=8'b11011110;
        13'd3376: m_out<=8'b11111001;
        13'd3377: m_out<=8'b11111111;
        13'd3378: m_out<=8'b11111101;
        13'd3379: m_out<=8'b11111110;
        13'd3380: m_out<=8'b11111110;
        13'd3381: m_out<=8'b11101011;
        13'd3382: m_out<=8'b11111000;
        13'd3383: m_out<=8'b11101010;
        13'd3384: m_out<=8'b00000110;
        13'd3385: m_out<=8'b11111000;
        13'd3386: m_out<=8'b11101110;
        13'd3387: m_out<=8'b00000010;
        13'd3388: m_out<=8'b11100000;
        13'd3389: m_out<=8'b00001111;
        13'd3390: m_out<=8'b00000011;
        13'd3391: m_out<=8'b00011000;
        13'd3392: m_out<=8'b11101000;
        13'd3393: m_out<=8'b11101111;
        13'd3394: m_out<=8'b00000011;
        13'd3395: m_out<=8'b00001101;
        13'd3396: m_out<=8'b00001110;
        13'd3397: m_out<=8'b11101001;
        13'd3398: m_out<=8'b11001000;
        13'd3399: m_out<=8'b11111010;
        13'd3400: m_out<=8'b00001110;
        13'd3401: m_out<=8'b11111000;
        13'd3402: m_out<=8'b11101110;
        13'd3403: m_out<=8'b11111110;
        13'd3404: m_out<=8'b11010111;
        13'd3405: m_out<=8'b00001011;
        13'd3406: m_out<=8'b11101010;
        13'd3407: m_out<=8'b00011000;
        13'd3408: m_out<=8'b11101011;
        13'd3409: m_out<=8'b00000001;
        13'd3410: m_out<=8'b00000111;
        13'd3411: m_out<=8'b00100111;
        13'd3412: m_out<=8'b11011011;
        13'd3413: m_out<=8'b00000010;
        13'd3414: m_out<=8'b11100100;
        13'd3415: m_out<=8'b00010101;
        13'd3416: m_out<=8'b11110111;
        13'd3417: m_out<=8'b11100001;
        13'd3418: m_out<=8'b00011111;
        13'd3419: m_out<=8'b00100010;
        13'd3420: m_out<=8'b11111000;
        13'd3421: m_out<=8'b11100000;
        13'd3422: m_out<=8'b11110011;
        13'd3423: m_out<=8'b00100110;
        13'd3424: m_out<=8'b11100000;
        13'd3425: m_out<=8'b00110001;
        13'd3426: m_out<=8'b00000011;
        13'd3427: m_out<=8'b11011100;
        13'd3428: m_out<=8'b00001110;
        13'd3429: m_out<=8'b11111100;
        13'd3430: m_out<=8'b00101011;
        13'd3431: m_out<=8'b11100001;
        13'd3432: m_out<=8'b11010101;
        13'd3433: m_out<=8'b11101110;
        13'd3434: m_out<=8'b00010110;
        13'd3435: m_out<=8'b11101000;
        13'd3436: m_out<=8'b11110111;
        13'd3437: m_out<=8'b11111100;
        13'd3438: m_out<=8'b11010100;
        13'd3439: m_out<=8'b11011010;
        13'd3440: m_out<=8'b00000111;
        13'd3441: m_out<=8'b00010001;
        13'd3442: m_out<=8'b11111101;
        13'd3443: m_out<=8'b11100100;
        13'd3444: m_out<=8'b00000111;
        13'd3445: m_out<=8'b00101000;
        13'd3446: m_out<=8'b00011100;
        13'd3447: m_out<=8'b11111001;
        13'd3448: m_out<=8'b11011010;
        13'd3449: m_out<=8'b01011011;
        13'd3450: m_out<=8'b00101010;
        13'd3451: m_out<=8'b11101000;
        13'd3452: m_out<=8'b00100110;
        13'd3453: m_out<=8'b11101011;
        13'd3454: m_out<=8'b11111100;
        13'd3455: m_out<=8'b11101101;
        13'd3456: m_out<=8'b00100010;
        13'd3457: m_out<=8'b11111001;
        13'd3458: m_out<=8'b00100000;
        13'd3459: m_out<=8'b00001010;
        13'd3460: m_out<=8'b00001100;
        13'd3461: m_out<=8'b11110110;
        13'd3462: m_out<=8'b00000111;
        13'd3463: m_out<=8'b00100011;
        13'd3464: m_out<=8'b11111011;
        13'd3465: m_out<=8'b11010000;
        13'd3466: m_out<=8'b11110101;
        13'd3467: m_out<=8'b11110001;
        13'd3468: m_out<=8'b10111100;
        13'd3469: m_out<=8'b00110000;
        13'd3470: m_out<=8'b11100000;
        13'd3471: m_out<=8'b11010011;
        13'd3472: m_out<=8'b00000110;
        13'd3473: m_out<=8'b11111001;
        13'd3474: m_out<=8'b11111011;
        13'd3475: m_out<=8'b11101100;
        13'd3476: m_out<=8'b00010101;
        13'd3477: m_out<=8'b11110111;
        13'd3478: m_out<=8'b11111011;
        13'd3479: m_out<=8'b00100100;
        13'd3480: m_out<=8'b00000101;
        13'd3481: m_out<=8'b00011100;
        13'd3482: m_out<=8'b00000011;
        13'd3483: m_out<=8'b00000101;
        13'd3484: m_out<=8'b11110100;
        13'd3485: m_out<=8'b00000001;
        13'd3486: m_out<=8'b00100010;
        13'd3487: m_out<=8'b00011011;
        13'd3488: m_out<=8'b00001110;
        13'd3489: m_out<=8'b00101111;
        13'd3490: m_out<=8'b00011100;
        13'd3491: m_out<=8'b00011111;
        13'd3492: m_out<=8'b00100101;
        13'd3493: m_out<=8'b00000001;
        13'd3494: m_out<=8'b11111010;
        13'd3495: m_out<=8'b00000000;
        13'd3496: m_out<=8'b00001110;
        13'd3497: m_out<=8'b11100110;
        13'd3498: m_out<=8'b11111000;
        13'd3499: m_out<=8'b11111100;
        13'd3500: m_out<=8'b00001011;
        13'd3501: m_out<=8'b00000000;
        13'd3502: m_out<=8'b11010001;
        13'd3503: m_out<=8'b00000110;
        13'd3504: m_out<=8'b11111000;
        13'd3505: m_out<=8'b00000101;
        13'd3506: m_out<=8'b00000100;
        13'd3507: m_out<=8'b11111110;
        13'd3508: m_out<=8'b11111100;
        13'd3509: m_out<=8'b11111110;
        13'd3510: m_out<=8'b00000011;
        13'd3511: m_out<=8'b11010011;
        13'd3512: m_out<=8'b00001000;
        13'd3513: m_out<=8'b00000111;
        13'd3514: m_out<=8'b11111110;
        13'd3515: m_out<=8'b00101111;
        13'd3516: m_out<=8'b11101111;
        13'd3517: m_out<=8'b00010101;
        13'd3518: m_out<=8'b11011010;
        13'd3519: m_out<=8'b11011001;
        13'd3520: m_out<=8'b00001000;
        13'd3521: m_out<=8'b00001011;
        13'd3522: m_out<=8'b00111011;
        13'd3523: m_out<=8'b00100001;
        13'd3524: m_out<=8'b11101000;
        13'd3525: m_out<=8'b00000110;
        13'd3526: m_out<=8'b00010001;
        13'd3527: m_out<=8'b00000101;
        13'd3528: m_out<=8'b11110111;
        13'd3529: m_out<=8'b11101000;
        13'd3530: m_out<=8'b11101110;
        13'd3531: m_out<=8'b00001101;
        13'd3532: m_out<=8'b11110001;
        13'd3533: m_out<=8'b00000000;
        13'd3534: m_out<=8'b11110000;
        13'd3535: m_out<=8'b11100110;
        13'd3536: m_out<=8'b11101101;
        13'd3537: m_out<=8'b00101101;
        13'd3538: m_out<=8'b00010100;
        13'd3539: m_out<=8'b00000001;
        13'd3540: m_out<=8'b00001000;
        13'd3541: m_out<=8'b11111101;
        13'd3542: m_out<=8'b00001001;
        13'd3543: m_out<=8'b00001001;
        13'd3544: m_out<=8'b00010010;
        13'd3545: m_out<=8'b00100000;
        13'd3546: m_out<=8'b00001101;
        13'd3547: m_out<=8'b11110010;
        13'd3548: m_out<=8'b11011100;
        13'd3549: m_out<=8'b00000001;
        13'd3550: m_out<=8'b11001100;
        13'd3551: m_out<=8'b11110100;
        13'd3552: m_out<=8'b11100001;
        13'd3553: m_out<=8'b00001011;
        13'd3554: m_out<=8'b11110101;
        13'd3555: m_out<=8'b11110000;
        13'd3556: m_out<=8'b11010110;
        13'd3557: m_out<=8'b11000111;
        13'd3558: m_out<=8'b11111100;
        13'd3559: m_out<=8'b00011010;
        13'd3560: m_out<=8'b00011100;
        13'd3561: m_out<=8'b11111110;
        13'd3562: m_out<=8'b11101000;
        13'd3563: m_out<=8'b11110110;
        13'd3564: m_out<=8'b00000001;
        13'd3565: m_out<=8'b11100011;
        13'd3566: m_out<=8'b11101110;
        13'd3567: m_out<=8'b00011010;
        13'd3568: m_out<=8'b00001111;
        13'd3569: m_out<=8'b11110010;
        13'd3570: m_out<=8'b11110011;
        13'd3571: m_out<=8'b11100100;
        13'd3572: m_out<=8'b11110010;
        13'd3573: m_out<=8'b00001111;
        13'd3574: m_out<=8'b11010100;
        13'd3575: m_out<=8'b11111011;
        13'd3576: m_out<=8'b00100000;
        13'd3577: m_out<=8'b11111101;
        13'd3578: m_out<=8'b11110100;
        13'd3579: m_out<=8'b00010001;
        13'd3580: m_out<=8'b00101000;
        13'd3581: m_out<=8'b11100000;
        13'd3582: m_out<=8'b00100001;
        13'd3583: m_out<=8'b11001110;
        13'd3584: m_out<=8'b11010010;
        13'd3585: m_out<=8'b00011101;
        13'd3586: m_out<=8'b11101110;
        13'd3587: m_out<=8'b00100000;
        13'd3588: m_out<=8'b11011110;
        13'd3589: m_out<=8'b11111100;
        13'd3590: m_out<=8'b00101000;
        13'd3591: m_out<=8'b00001010;
        13'd3592: m_out<=8'b00001110;
        13'd3593: m_out<=8'b00000011;
        13'd3594: m_out<=8'b00000110;
        13'd3595: m_out<=8'b11111111;
        13'd3596: m_out<=8'b11011100;
        13'd3597: m_out<=8'b11111101;
        13'd3598: m_out<=8'b00000000;
        13'd3599: m_out<=8'b00101010;
        13'd3600: m_out<=8'b00000101;
        13'd3601: m_out<=8'b11101101;
        13'd3602: m_out<=8'b00011000;
        13'd3603: m_out<=8'b00001100;
        13'd3604: m_out<=8'b11000101;
        13'd3605: m_out<=8'b11010101;
        13'd3606: m_out<=8'b00100100;
        13'd3607: m_out<=8'b00110111;
        13'd3608: m_out<=8'b00000011;
        13'd3609: m_out<=8'b11011001;
        13'd3610: m_out<=8'b11100110;
        13'd3611: m_out<=8'b00001100;
        13'd3612: m_out<=8'b11011000;
        13'd3613: m_out<=8'b00000100;
        13'd3614: m_out<=8'b00010101;
        13'd3615: m_out<=8'b11110110;
        13'd3616: m_out<=8'b01000010;
        13'd3617: m_out<=8'b00010101;
        13'd3618: m_out<=8'b00100010;
        13'd3619: m_out<=8'b00001110;
        13'd3620: m_out<=8'b11101100;
        13'd3621: m_out<=8'b11100011;
        13'd3622: m_out<=8'b00000011;
        13'd3623: m_out<=8'b00100011;
        13'd3624: m_out<=8'b00000100;
        13'd3625: m_out<=8'b00000111;
        13'd3626: m_out<=8'b00100011;
        13'd3627: m_out<=8'b00101100;
        13'd3628: m_out<=8'b00000101;
        13'd3629: m_out<=8'b00010001;
        13'd3630: m_out<=8'b11110000;
        13'd3631: m_out<=8'b11100001;
        13'd3632: m_out<=8'b00011010;
        13'd3633: m_out<=8'b11111011;
        13'd3634: m_out<=8'b00000100;
        13'd3635: m_out<=8'b11101101;
        13'd3636: m_out<=8'b11101010;
        13'd3637: m_out<=8'b00011101;
        13'd3638: m_out<=8'b11100010;
        13'd3639: m_out<=8'b11100011;
        13'd3640: m_out<=8'b00011110;
        13'd3641: m_out<=8'b11110011;
        13'd3642: m_out<=8'b11111100;
        13'd3643: m_out<=8'b00100111;
        13'd3644: m_out<=8'b11111010;
        13'd3645: m_out<=8'b11111111;
        13'd3646: m_out<=8'b11101100;
        13'd3647: m_out<=8'b11000110;
        13'd3648: m_out<=8'b00011011;
        13'd3649: m_out<=8'b00100101;
        13'd3650: m_out<=8'b11011111;
        13'd3651: m_out<=8'b11010101;
        13'd3652: m_out<=8'b00001101;
        13'd3653: m_out<=8'b11101100;
        13'd3654: m_out<=8'b11101101;
        13'd3655: m_out<=8'b11001001;
        13'd3656: m_out<=8'b00001111;
        13'd3657: m_out<=8'b11101101;
        13'd3658: m_out<=8'b00010011;
        13'd3659: m_out<=8'b11100101;
        13'd3660: m_out<=8'b00000111;
        13'd3661: m_out<=8'b00011111;
        13'd3662: m_out<=8'b10111100;
        13'd3663: m_out<=8'b00000101;
        13'd3664: m_out<=8'b11110000;
        13'd3665: m_out<=8'b00100111;
        13'd3666: m_out<=8'b11110110;
        13'd3667: m_out<=8'b00000110;
        13'd3668: m_out<=8'b00010111;
        13'd3669: m_out<=8'b00000001;
        13'd3670: m_out<=8'b00000110;
        13'd3671: m_out<=8'b00010001;
        13'd3672: m_out<=8'b11110000;
        13'd3673: m_out<=8'b00010111;
        13'd3674: m_out<=8'b00010000;
        13'd3675: m_out<=8'b00011110;
        13'd3676: m_out<=8'b11111111;
        13'd3677: m_out<=8'b11110001;
        13'd3678: m_out<=8'b00000110;
        13'd3679: m_out<=8'b00000000;
        13'd3680: m_out<=8'b00010100;
        13'd3681: m_out<=8'b00010010;
        13'd3682: m_out<=8'b11101010;
        13'd3683: m_out<=8'b00010100;
        13'd3684: m_out<=8'b11101111;
        13'd3685: m_out<=8'b00000001;
        13'd3686: m_out<=8'b00010011;
        13'd3687: m_out<=8'b00011000;
        13'd3688: m_out<=8'b01001000;
        13'd3689: m_out<=8'b00010011;
        13'd3690: m_out<=8'b11010111;
        13'd3691: m_out<=8'b11101001;
        13'd3692: m_out<=8'b00001100;
        13'd3693: m_out<=8'b00000111;
        13'd3694: m_out<=8'b00010101;
        13'd3695: m_out<=8'b00100100;
        13'd3696: m_out<=8'b00000001;
        13'd3697: m_out<=8'b00001110;
        13'd3698: m_out<=8'b11111111;
        13'd3699: m_out<=8'b11101101;
        13'd3700: m_out<=8'b00011000;
        13'd3701: m_out<=8'b11111001;
        13'd3702: m_out<=8'b11111100;
        13'd3703: m_out<=8'b11110001;
        13'd3704: m_out<=8'b11111101;
        13'd3705: m_out<=8'b00000010;
        13'd3706: m_out<=8'b11101111;
        13'd3707: m_out<=8'b11101110;
        13'd3708: m_out<=8'b11110011;
        13'd3709: m_out<=8'b00010011;
        13'd3710: m_out<=8'b11101111;
        13'd3711: m_out<=8'b00000111;
        13'd3712: m_out<=8'b11110110;
        13'd3713: m_out<=8'b00000110;
        13'd3714: m_out<=8'b00001101;
        13'd3715: m_out<=8'b00001001;
        13'd3716: m_out<=8'b00000001;
        13'd3717: m_out<=8'b11101100;
        13'd3718: m_out<=8'b00101110;
        13'd3719: m_out<=8'b00100100;
        13'd3720: m_out<=8'b11101100;
        13'd3721: m_out<=8'b00000011;
        13'd3722: m_out<=8'b00001110;
        13'd3723: m_out<=8'b11011011;
        13'd3724: m_out<=8'b11111011;
        13'd3725: m_out<=8'b00010001;
        13'd3726: m_out<=8'b11100101;
        13'd3727: m_out<=8'b11100101;
        13'd3728: m_out<=8'b00011011;
        13'd3729: m_out<=8'b11101101;
        13'd3730: m_out<=8'b11111001;
        13'd3731: m_out<=8'b00110100;
        13'd3732: m_out<=8'b00110000;
        13'd3733: m_out<=8'b11101011;
        13'd3734: m_out<=8'b00101010;
        13'd3735: m_out<=8'b11101111;
        13'd3736: m_out<=8'b11000100;
        13'd3737: m_out<=8'b11111011;
        13'd3738: m_out<=8'b11111000;
        13'd3739: m_out<=8'b11110001;
        13'd3740: m_out<=8'b00001010;
        13'd3741: m_out<=8'b11100101;
        13'd3742: m_out<=8'b11010100;
        13'd3743: m_out<=8'b00101001;
        13'd3744: m_out<=8'b00101000;
        13'd3745: m_out<=8'b00001111;
        13'd3746: m_out<=8'b00010011;
        13'd3747: m_out<=8'b00001100;
        13'd3748: m_out<=8'b00100111;
        13'd3749: m_out<=8'b00101000;
        13'd3750: m_out<=8'b11100001;
        13'd3751: m_out<=8'b11110001;
        13'd3752: m_out<=8'b00001000;
        13'd3753: m_out<=8'b00110100;
        13'd3754: m_out<=8'b11101011;
        13'd3755: m_out<=8'b01011010;
        13'd3756: m_out<=8'b11110110;
        13'd3757: m_out<=8'b11110110;
        13'd3758: m_out<=8'b11100000;
        13'd3759: m_out<=8'b00000101;
        13'd3760: m_out<=8'b00100010;
        13'd3761: m_out<=8'b00010001;
        13'd3762: m_out<=8'b00010100;
        13'd3763: m_out<=8'b11100101;
        13'd3764: m_out<=8'b11100001;
        13'd3765: m_out<=8'b00000000;
        13'd3766: m_out<=8'b11111101;
        13'd3767: m_out<=8'b11111001;
        13'd3768: m_out<=8'b00010001;
        13'd3769: m_out<=8'b11111010;
        13'd3770: m_out<=8'b00101001;
        13'd3771: m_out<=8'b00000100;
        13'd3772: m_out<=8'b11110101;
        13'd3773: m_out<=8'b00010001;
        13'd3774: m_out<=8'b00001111;
        13'd3775: m_out<=8'b00000100;
        13'd3776: m_out<=8'b00000000;
        13'd3777: m_out<=8'b00000111;
        13'd3778: m_out<=8'b00101101;
        13'd3779: m_out<=8'b00000100;
        13'd3780: m_out<=8'b00001010;
        13'd3781: m_out<=8'b00000110;
        13'd3782: m_out<=8'b11101000;
        13'd3783: m_out<=8'b00010001;
        13'd3784: m_out<=8'b11110010;
        13'd3785: m_out<=8'b11100111;
        13'd3786: m_out<=8'b00010010;
        13'd3787: m_out<=8'b11111111;
        13'd3788: m_out<=8'b00000010;
        13'd3789: m_out<=8'b11010001;
        13'd3790: m_out<=8'b11111010;
        13'd3791: m_out<=8'b00000100;
        13'd3792: m_out<=8'b11111110;
        13'd3793: m_out<=8'b00001011;
        13'd3794: m_out<=8'b00111100;
        13'd3795: m_out<=8'b00100110;
        13'd3796: m_out<=8'b11111111;
        13'd3797: m_out<=8'b11110111;
        13'd3798: m_out<=8'b00011011;
        13'd3799: m_out<=8'b00000111;
        13'd3800: m_out<=8'b11110011;
        13'd3801: m_out<=8'b11111101;
        13'd3802: m_out<=8'b11101100;
        13'd3803: m_out<=8'b11100101;
        13'd3804: m_out<=8'b00010101;
        13'd3805: m_out<=8'b00001011;
        13'd3806: m_out<=8'b00011111;
        13'd3807: m_out<=8'b11101011;
        13'd3808: m_out<=8'b00000010;
        13'd3809: m_out<=8'b11111000;
        13'd3810: m_out<=8'b00001010;
        13'd3811: m_out<=8'b00000011;
        13'd3812: m_out<=8'b11110101;
        13'd3813: m_out<=8'b00110110;
        13'd3814: m_out<=8'b11111100;
        13'd3815: m_out<=8'b00011100;
        13'd3816: m_out<=8'b00001100;
        13'd3817: m_out<=8'b11010111;
        13'd3818: m_out<=8'b00001101;
        13'd3819: m_out<=8'b11111101;
        13'd3820: m_out<=8'b00011110;
        13'd3821: m_out<=8'b00011000;
        13'd3822: m_out<=8'b00000010;
        13'd3823: m_out<=8'b11010110;
        13'd3824: m_out<=8'b00011010;
        13'd3825: m_out<=8'b00010110;
        13'd3826: m_out<=8'b00011010;
        13'd3827: m_out<=8'b11101110;
        13'd3828: m_out<=8'b00000001;
        13'd3829: m_out<=8'b00100100;
        13'd3830: m_out<=8'b00001010;
        13'd3831: m_out<=8'b00000101;
        13'd3832: m_out<=8'b11111010;
        13'd3833: m_out<=8'b11110011;
        13'd3834: m_out<=8'b00101101;
        13'd3835: m_out<=8'b00001001;
        13'd3836: m_out<=8'b11100010;
        13'd3837: m_out<=8'b00000000;
        13'd3838: m_out<=8'b11110100;
        13'd3839: m_out<=8'b11101100;
        13'd3840: m_out<=8'b10101110;
        13'd3841: m_out<=8'b00000110;
        13'd3842: m_out<=8'b00000101;
        13'd3843: m_out<=8'b00001101;
        13'd3844: m_out<=8'b11110100;
        13'd3845: m_out<=8'b11010110;
        13'd3846: m_out<=8'b00001011;
        13'd3847: m_out<=8'b11110000;
        13'd3848: m_out<=8'b00011011;
        13'd3849: m_out<=8'b00000111;
        13'd3850: m_out<=8'b11110111;
        13'd3851: m_out<=8'b00110001;
        13'd3852: m_out<=8'b00011100;
        13'd3853: m_out<=8'b11110011;
        13'd3854: m_out<=8'b00010110;
        13'd3855: m_out<=8'b11011110;
        13'd3856: m_out<=8'b00111011;
        13'd3857: m_out<=8'b11011110;
        13'd3858: m_out<=8'b00010111;
        13'd3859: m_out<=8'b11110111;
        13'd3860: m_out<=8'b11101010;
        13'd3861: m_out<=8'b00010111;
        13'd3862: m_out<=8'b00011100;
        13'd3863: m_out<=8'b11101101;
        13'd3864: m_out<=8'b11110000;
        13'd3865: m_out<=8'b00000100;
        13'd3866: m_out<=8'b11110011;
        13'd3867: m_out<=8'b00010011;
        13'd3868: m_out<=8'b10111101;
        13'd3869: m_out<=8'b00000100;
        13'd3870: m_out<=8'b00000110;
        13'd3871: m_out<=8'b11011011;
        13'd3872: m_out<=8'b00001001;
        13'd3873: m_out<=8'b11111010;
        13'd3874: m_out<=8'b11111111;
        13'd3875: m_out<=8'b11111111;
        13'd3876: m_out<=8'b11110001;
        13'd3877: m_out<=8'b00100101;
        13'd3878: m_out<=8'b11001101;
        13'd3879: m_out<=8'b11101111;
        13'd3880: m_out<=8'b11000100;
        13'd3881: m_out<=8'b00011011;
        13'd3882: m_out<=8'b11100110;
        13'd3883: m_out<=8'b00011011;
        13'd3884: m_out<=8'b00001100;
        13'd3885: m_out<=8'b00110110;
        13'd3886: m_out<=8'b00000110;
        13'd3887: m_out<=8'b11111100;
        13'd3888: m_out<=8'b11110101;
        13'd3889: m_out<=8'b00011100;
        13'd3890: m_out<=8'b11011101;
        13'd3891: m_out<=8'b00001001;
        13'd3892: m_out<=8'b00101101;
        13'd3893: m_out<=8'b11101101;
        13'd3894: m_out<=8'b00000010;
        13'd3895: m_out<=8'b00000010;
        13'd3896: m_out<=8'b11101010;
        13'd3897: m_out<=8'b11101100;
        13'd3898: m_out<=8'b00000110;
        13'd3899: m_out<=8'b11101110;
        13'd3900: m_out<=8'b11110011;
        13'd3901: m_out<=8'b11110110;
        13'd3902: m_out<=8'b11110110;
        13'd3903: m_out<=8'b00001101;
        13'd3904: m_out<=8'b11111010;
        13'd3905: m_out<=8'b00100100;
        13'd3906: m_out<=8'b00010010;
        13'd3907: m_out<=8'b11101100;
        13'd3908: m_out<=8'b00000010;
        13'd3909: m_out<=8'b00000110;
        13'd3910: m_out<=8'b00110111;
        13'd3911: m_out<=8'b11110111;
        13'd3912: m_out<=8'b00100100;
        13'd3913: m_out<=8'b00010100;
        13'd3914: m_out<=8'b00100000;
        13'd3915: m_out<=8'b00000000;
        13'd3916: m_out<=8'b11111011;
        13'd3917: m_out<=8'b11100111;
        13'd3918: m_out<=8'b00001100;
        13'd3919: m_out<=8'b11101101;
        13'd3920: m_out<=8'b11111111;
        13'd3921: m_out<=8'b00000111;
        13'd3922: m_out<=8'b00001011;
        13'd3923: m_out<=8'b11001010;
        13'd3924: m_out<=8'b11010010;
        13'd3925: m_out<=8'b00110000;
        13'd3926: m_out<=8'b11010010;
        13'd3927: m_out<=8'b00010011;
        13'd3928: m_out<=8'b11001110;
        13'd3929: m_out<=8'b11101111;
        13'd3930: m_out<=8'b11111110;
        13'd3931: m_out<=8'b11101010;
        13'd3932: m_out<=8'b11010110;
        13'd3933: m_out<=8'b00010010;
        13'd3934: m_out<=8'b11100100;
        13'd3935: m_out<=8'b11101100;
        13'd3936: m_out<=8'b00000000;
        13'd3937: m_out<=8'b11110100;
        13'd3938: m_out<=8'b00001110;
        13'd3939: m_out<=8'b11111001;
        13'd3940: m_out<=8'b00011100;
        13'd3941: m_out<=8'b11010000;
        13'd3942: m_out<=8'b11111110;
        13'd3943: m_out<=8'b11110001;
        13'd3944: m_out<=8'b11100011;
        13'd3945: m_out<=8'b00100001;
        13'd3946: m_out<=8'b00000001;
        13'd3947: m_out<=8'b11110010;
        13'd3948: m_out<=8'b11111101;
        13'd3949: m_out<=8'b00110111;
        13'd3950: m_out<=8'b11110010;
        13'd3951: m_out<=8'b11011100;
        13'd3952: m_out<=8'b00100101;
        13'd3953: m_out<=8'b11110011;
        13'd3954: m_out<=8'b00010000;
        13'd3955: m_out<=8'b00011000;
        13'd3956: m_out<=8'b00001000;
        13'd3957: m_out<=8'b00011011;
        13'd3958: m_out<=8'b11110001;
        13'd3959: m_out<=8'b00100001;
        13'd3960: m_out<=8'b11001100;
        13'd3961: m_out<=8'b00101100;
        13'd3962: m_out<=8'b11011011;
        13'd3963: m_out<=8'b11000001;
        13'd3964: m_out<=8'b00000111;
        13'd3965: m_out<=8'b00000101;
        13'd3966: m_out<=8'b11100101;
        13'd3967: m_out<=8'b11101110;
        13'd3968: m_out<=8'b00100001;
        13'd3969: m_out<=8'b00011001;
        13'd3970: m_out<=8'b00010110;
        13'd3971: m_out<=8'b11101010;
        13'd3972: m_out<=8'b11110101;
        13'd3973: m_out<=8'b00011111;
        13'd3974: m_out<=8'b11111011;
        13'd3975: m_out<=8'b11110011;
        13'd3976: m_out<=8'b11111110;
        13'd3977: m_out<=8'b00011001;
        13'd3978: m_out<=8'b11011111;
        13'd3979: m_out<=8'b11100001;
        13'd3980: m_out<=8'b00001111;
        13'd3981: m_out<=8'b00010111;
        13'd3982: m_out<=8'b00000100;
        13'd3983: m_out<=8'b00010101;
        13'd3984: m_out<=8'b11110001;
        13'd3985: m_out<=8'b00010011;
        13'd3986: m_out<=8'b11010101;
        13'd3987: m_out<=8'b00011101;
        13'd3988: m_out<=8'b00101101;
        13'd3989: m_out<=8'b00000000;
        13'd3990: m_out<=8'b00010001;
        13'd3991: m_out<=8'b00001001;
        13'd3992: m_out<=8'b00010000;
        13'd3993: m_out<=8'b00001101;
        13'd3994: m_out<=8'b11110000;
        13'd3995: m_out<=8'b00001101;
        13'd3996: m_out<=8'b00001100;
        13'd3997: m_out<=8'b11101110;
        13'd3998: m_out<=8'b11101000;
        13'd3999: m_out<=8'b11111111;
        13'd4000: m_out<=8'b00001101;
        13'd4001: m_out<=8'b11111010;
        13'd4002: m_out<=8'b11111011;
        13'd4003: m_out<=8'b00010000;
        13'd4004: m_out<=8'b00011000;
        13'd4005: m_out<=8'b00010111;
        13'd4006: m_out<=8'b11100110;
        13'd4007: m_out<=8'b11011010;
        13'd4008: m_out<=8'b11110010;
        13'd4009: m_out<=8'b00001100;
        13'd4010: m_out<=8'b11110111;
        13'd4011: m_out<=8'b00000111;
        13'd4012: m_out<=8'b00010110;
        13'd4013: m_out<=8'b00001011;
        13'd4014: m_out<=8'b00000110;
        13'd4015: m_out<=8'b00010011;
        13'd4016: m_out<=8'b11100110;
        13'd4017: m_out<=8'b00011001;
        13'd4018: m_out<=8'b00011000;
        13'd4019: m_out<=8'b00110001;
        13'd4020: m_out<=8'b00000110;
        13'd4021: m_out<=8'b00001101;
        13'd4022: m_out<=8'b11100100;
        13'd4023: m_out<=8'b00011000;
        13'd4024: m_out<=8'b11110111;
        13'd4025: m_out<=8'b00011001;
        13'd4026: m_out<=8'b00000011;
        13'd4027: m_out<=8'b11111110;
        13'd4028: m_out<=8'b00001111;
        13'd4029: m_out<=8'b00000011;
        13'd4030: m_out<=8'b00100010;
        13'd4031: m_out<=8'b00101000;
        13'd4032: m_out<=8'b00100000;
        13'd4033: m_out<=8'b11110010;
        13'd4034: m_out<=8'b11110101;
        13'd4035: m_out<=8'b11111000;
        13'd4036: m_out<=8'b00010110;
        13'd4037: m_out<=8'b00001110;
        13'd4038: m_out<=8'b00001000;
        13'd4039: m_out<=8'b11001011;
        13'd4040: m_out<=8'b11010110;
        13'd4041: m_out<=8'b00000000;
        13'd4042: m_out<=8'b11101111;
        13'd4043: m_out<=8'b00010100;
        13'd4044: m_out<=8'b00000001;
        13'd4045: m_out<=8'b00110011;
        13'd4046: m_out<=8'b00001101;
        13'd4047: m_out<=8'b11100101;
        13'd4048: m_out<=8'b11110110;
        13'd4049: m_out<=8'b11110111;
        13'd4050: m_out<=8'b00001101;
        13'd4051: m_out<=8'b00000110;
        13'd4052: m_out<=8'b11101000;
        13'd4053: m_out<=8'b11111011;
        13'd4054: m_out<=8'b11111000;
        13'd4055: m_out<=8'b00010110;
        13'd4056: m_out<=8'b00001000;
        13'd4057: m_out<=8'b11110000;
        13'd4058: m_out<=8'b00000011;
        13'd4059: m_out<=8'b00001001;
        13'd4060: m_out<=8'b11011100;
        13'd4061: m_out<=8'b11111001;
        13'd4062: m_out<=8'b00010000;
        13'd4063: m_out<=8'b00000101;
        13'd4064: m_out<=8'b00010000;
        13'd4065: m_out<=8'b00011010;
        13'd4066: m_out<=8'b11111010;
        13'd4067: m_out<=8'b00001101;
        13'd4068: m_out<=8'b00000010;
        13'd4069: m_out<=8'b11101011;
        13'd4070: m_out<=8'b11100001;
        13'd4071: m_out<=8'b00000001;
        13'd4072: m_out<=8'b00100111;
        13'd4073: m_out<=8'b11011010;
        13'd4074: m_out<=8'b11111101;
        13'd4075: m_out<=8'b00000110;
        13'd4076: m_out<=8'b11001100;
        13'd4077: m_out<=8'b00010111;
        13'd4078: m_out<=8'b11111000;
        13'd4079: m_out<=8'b00000110;
        13'd4080: m_out<=8'b00001110;
        13'd4081: m_out<=8'b11110000;
        13'd4082: m_out<=8'b00101010;
        13'd4083: m_out<=8'b00001101;
        13'd4084: m_out<=8'b00011111;
        13'd4085: m_out<=8'b00001100;
        13'd4086: m_out<=8'b11110111;
        13'd4087: m_out<=8'b11101011;
        13'd4088: m_out<=8'b11011110;
        13'd4089: m_out<=8'b00000100;
        13'd4090: m_out<=8'b00000100;
        13'd4091: m_out<=8'b00001110;
        13'd4092: m_out<=8'b00011001;
        13'd4093: m_out<=8'b00010011;
        13'd4094: m_out<=8'b00100110;
        13'd4095: m_out<=8'b11010100;
        13'd4096: m_out<=8'b00001100;
        13'd4097: m_out<=8'b00011100;
        13'd4098: m_out<=8'b00001111;
        13'd4099: m_out<=8'b11111011;
        13'd4100: m_out<=8'b11011110;
        13'd4101: m_out<=8'b00010010;
        13'd4102: m_out<=8'b11100011;
        13'd4103: m_out<=8'b11110101;
        13'd4104: m_out<=8'b11110110;
        13'd4105: m_out<=8'b11100001;
        13'd4106: m_out<=8'b00000100;
        13'd4107: m_out<=8'b00011001;
        13'd4108: m_out<=8'b00011100;
        13'd4109: m_out<=8'b00000100;
        13'd4110: m_out<=8'b00110110;
        13'd4111: m_out<=8'b00010011;
        13'd4112: m_out<=8'b00001101;
        13'd4113: m_out<=8'b11111001;
        13'd4114: m_out<=8'b00000111;
        13'd4115: m_out<=8'b11100001;
        13'd4116: m_out<=8'b00011001;
        13'd4117: m_out<=8'b00010101;
        13'd4118: m_out<=8'b11110111;
        13'd4119: m_out<=8'b11010000;
        13'd4120: m_out<=8'b11101010;
        13'd4121: m_out<=8'b00000110;
        13'd4122: m_out<=8'b11110000;
        13'd4123: m_out<=8'b11010111;
        13'd4124: m_out<=8'b11011001;
        13'd4125: m_out<=8'b00010011;
        13'd4126: m_out<=8'b00011001;
        13'd4127: m_out<=8'b00001101;
        13'd4128: m_out<=8'b00000110;
        13'd4129: m_out<=8'b11111001;
        13'd4130: m_out<=8'b11101000;
        13'd4131: m_out<=8'b11101011;
        13'd4132: m_out<=8'b00000000;
        13'd4133: m_out<=8'b00001000;
        13'd4134: m_out<=8'b00001011;
        13'd4135: m_out<=8'b11111101;
        13'd4136: m_out<=8'b00001001;
        13'd4137: m_out<=8'b00101011;
        13'd4138: m_out<=8'b00010101;
        13'd4139: m_out<=8'b00100011;
        13'd4140: m_out<=8'b00100110;
        13'd4141: m_out<=8'b11101111;
        13'd4142: m_out<=8'b00111101;
        13'd4143: m_out<=8'b00011000;
        13'd4144: m_out<=8'b11111011;
        13'd4145: m_out<=8'b00000011;
        13'd4146: m_out<=8'b11111100;
        13'd4147: m_out<=8'b00100001;
        13'd4148: m_out<=8'b00011000;
        13'd4149: m_out<=8'b00001100;
        13'd4150: m_out<=8'b11101010;
        13'd4151: m_out<=8'b00100101;
        13'd4152: m_out<=8'b00101001;
        13'd4153: m_out<=8'b00101000;
        13'd4154: m_out<=8'b11100111;
        13'd4155: m_out<=8'b00110001;
        13'd4156: m_out<=8'b00010010;
        13'd4157: m_out<=8'b00000010;
        13'd4158: m_out<=8'b00001010;
        13'd4159: m_out<=8'b00010100;
        13'd4160: m_out<=8'b11011100;
        13'd4161: m_out<=8'b00010101;
        13'd4162: m_out<=8'b00000100;
        13'd4163: m_out<=8'b00011010;
        13'd4164: m_out<=8'b00001100;
        13'd4165: m_out<=8'b11111100;
        13'd4166: m_out<=8'b00001110;
        13'd4167: m_out<=8'b11111111;
        13'd4168: m_out<=8'b00100001;
        13'd4169: m_out<=8'b11000101;
        13'd4170: m_out<=8'b11100110;
        13'd4171: m_out<=8'b11110111;
        13'd4172: m_out<=8'b11111100;
        13'd4173: m_out<=8'b00000011;
        13'd4174: m_out<=8'b00100010;
        13'd4175: m_out<=8'b00010101;
        13'd4176: m_out<=8'b11100111;
        13'd4177: m_out<=8'b00000010;
        13'd4178: m_out<=8'b00010101;
        13'd4179: m_out<=8'b11101011;
        13'd4180: m_out<=8'b11101001;
        13'd4181: m_out<=8'b00101111;
        13'd4182: m_out<=8'b00111110;
        13'd4183: m_out<=8'b11100101;
        13'd4184: m_out<=8'b00011000;
        13'd4185: m_out<=8'b00010111;
        13'd4186: m_out<=8'b11100001;
        13'd4187: m_out<=8'b11110111;
        13'd4188: m_out<=8'b11111111;
        13'd4189: m_out<=8'b00000001;
        13'd4190: m_out<=8'b11101011;
        13'd4191: m_out<=8'b11110000;
        13'd4192: m_out<=8'b00011010;
        13'd4193: m_out<=8'b00000010;
        13'd4194: m_out<=8'b11111001;
        13'd4195: m_out<=8'b11100001;
        13'd4196: m_out<=8'b00010110;
        13'd4197: m_out<=8'b11110001;
        13'd4198: m_out<=8'b11000011;
        13'd4199: m_out<=8'b11011001;
        13'd4200: m_out<=8'b11100110;
        13'd4201: m_out<=8'b11110001;
        13'd4202: m_out<=8'b11110000;
        13'd4203: m_out<=8'b00001111;
        13'd4204: m_out<=8'b00001001;
        13'd4205: m_out<=8'b11111111;
        13'd4206: m_out<=8'b11011101;
        13'd4207: m_out<=8'b00111010;
        13'd4208: m_out<=8'b00010100;
        13'd4209: m_out<=8'b00001000;
        13'd4210: m_out<=8'b11100011;
        13'd4211: m_out<=8'b11110010;
        13'd4212: m_out<=8'b00011000;
        13'd4213: m_out<=8'b00100011;
        13'd4214: m_out<=8'b11101111;
        13'd4215: m_out<=8'b11110010;
        13'd4216: m_out<=8'b00010110;
        13'd4217: m_out<=8'b00010110;
        13'd4218: m_out<=8'b00000011;
        13'd4219: m_out<=8'b00001110;
        13'd4220: m_out<=8'b00000100;
        13'd4221: m_out<=8'b00000001;
        13'd4222: m_out<=8'b11111110;
        13'd4223: m_out<=8'b00001101;
        13'd4224: m_out<=8'b11111101;
        13'd4225: m_out<=8'b11111111;
        13'd4226: m_out<=8'b00000100;
        13'd4227: m_out<=8'b11110101;
        13'd4228: m_out<=8'b11011111;
        13'd4229: m_out<=8'b11011110;
        13'd4230: m_out<=8'b00001000;
        13'd4231: m_out<=8'b00000000;
        13'd4232: m_out<=8'b00010001;
        13'd4233: m_out<=8'b11100011;
        13'd4234: m_out<=8'b00001100;
        13'd4235: m_out<=8'b11101010;
        13'd4236: m_out<=8'b00000001;
        13'd4237: m_out<=8'b11111110;
        13'd4238: m_out<=8'b00001110;
        13'd4239: m_out<=8'b00010011;
        13'd4240: m_out<=8'b00011110;
        13'd4241: m_out<=8'b00111110;
        13'd4242: m_out<=8'b00011010;
        13'd4243: m_out<=8'b00001000;
        13'd4244: m_out<=8'b00000111;
        13'd4245: m_out<=8'b00010011;
        13'd4246: m_out<=8'b11011010;
        13'd4247: m_out<=8'b11101001;
        13'd4248: m_out<=8'b11000111;
        13'd4249: m_out<=8'b00001101;
        13'd4250: m_out<=8'b11011111;
        13'd4251: m_out<=8'b11110111;
        13'd4252: m_out<=8'b11111100;
        13'd4253: m_out<=8'b00110101;
        13'd4254: m_out<=8'b11011000;
        13'd4255: m_out<=8'b00000000;
        13'd4256: m_out<=8'b00010100;
        13'd4257: m_out<=8'b00000001;
        13'd4258: m_out<=8'b00100011;
        13'd4259: m_out<=8'b00001001;
        13'd4260: m_out<=8'b00001101;
        13'd4261: m_out<=8'b11100000;
        13'd4262: m_out<=8'b11100110;
        13'd4263: m_out<=8'b00001100;
        13'd4264: m_out<=8'b00001101;
        13'd4265: m_out<=8'b11001001;
        13'd4266: m_out<=8'b00010110;
        13'd4267: m_out<=8'b11011000;
        13'd4268: m_out<=8'b11100100;
        13'd4269: m_out<=8'b00010011;
        13'd4270: m_out<=8'b00001111;
        13'd4271: m_out<=8'b11100011;
        13'd4272: m_out<=8'b00001011;
        13'd4273: m_out<=8'b00100100;
        13'd4274: m_out<=8'b00111111;
        13'd4275: m_out<=8'b11000101;
        13'd4276: m_out<=8'b11111110;
        13'd4277: m_out<=8'b11110000;
        13'd4278: m_out<=8'b00010001;
        13'd4279: m_out<=8'b11100100;
        13'd4280: m_out<=8'b00100110;
        13'd4281: m_out<=8'b11111111;
        13'd4282: m_out<=8'b00010001;
        13'd4283: m_out<=8'b00110100;
        13'd4284: m_out<=8'b11011010;
        13'd4285: m_out<=8'b00000110;
        13'd4286: m_out<=8'b11111110;
        13'd4287: m_out<=8'b00011010;
        13'd4288: m_out<=8'b11101001;
        13'd4289: m_out<=8'b11110111;
        13'd4290: m_out<=8'b00011110;
        13'd4291: m_out<=8'b00010001;
        13'd4292: m_out<=8'b00011110;
        13'd4293: m_out<=8'b00000011;
        13'd4294: m_out<=8'b00001010;
        13'd4295: m_out<=8'b00100001;
        13'd4296: m_out<=8'b11110101;
        13'd4297: m_out<=8'b00000111;
        13'd4298: m_out<=8'b00001110;
        13'd4299: m_out<=8'b11110110;
        13'd4300: m_out<=8'b11011111;
        13'd4301: m_out<=8'b11110111;
        13'd4302: m_out<=8'b00000101;
        13'd4303: m_out<=8'b00001011;
        13'd4304: m_out<=8'b11110110;
        13'd4305: m_out<=8'b00100101;
        13'd4306: m_out<=8'b11111010;
        13'd4307: m_out<=8'b00110100;
        13'd4308: m_out<=8'b00010010;
        13'd4309: m_out<=8'b00010010;
        13'd4310: m_out<=8'b11111100;
        13'd4311: m_out<=8'b11100101;
        13'd4312: m_out<=8'b00011010;
        13'd4313: m_out<=8'b00011110;
        13'd4314: m_out<=8'b11011011;
        13'd4315: m_out<=8'b00010111;
        13'd4316: m_out<=8'b11101100;
        13'd4317: m_out<=8'b00111001;
        13'd4318: m_out<=8'b00000111;
        13'd4319: m_out<=8'b00001111;
        13'd4320: m_out<=8'b10101101;
        13'd4321: m_out<=8'b11111100;
        13'd4322: m_out<=8'b00000000;
        13'd4323: m_out<=8'b11011000;
        13'd4324: m_out<=8'b11110111;
        13'd4325: m_out<=8'b00000011;
        13'd4326: m_out<=8'b00010001;
        13'd4327: m_out<=8'b00011010;
        13'd4328: m_out<=8'b11110100;
        13'd4329: m_out<=8'b11110001;
        13'd4330: m_out<=8'b00001110;
        13'd4331: m_out<=8'b00001100;
        13'd4332: m_out<=8'b00000100;
        13'd4333: m_out<=8'b11110100;
        13'd4334: m_out<=8'b00100000;
        13'd4335: m_out<=8'b00001010;
        13'd4336: m_out<=8'b00010000;
        13'd4337: m_out<=8'b00010001;
        13'd4338: m_out<=8'b00011110;
        13'd4339: m_out<=8'b00001110;
        13'd4340: m_out<=8'b00000010;
        13'd4341: m_out<=8'b00000011;
        13'd4342: m_out<=8'b11110100;
        13'd4343: m_out<=8'b00000100;
        13'd4344: m_out<=8'b00000111;
        13'd4345: m_out<=8'b00001000;
        13'd4346: m_out<=8'b00011100;
        13'd4347: m_out<=8'b01001001;
        13'd4348: m_out<=8'b00001011;
        13'd4349: m_out<=8'b11100000;
        13'd4350: m_out<=8'b11111011;
        13'd4351: m_out<=8'b00000000;
        13'd4352: m_out<=8'b11100100;
        13'd4353: m_out<=8'b11000110;
        13'd4354: m_out<=8'b00001110;
        13'd4355: m_out<=8'b00000000;
        13'd4356: m_out<=8'b11101111;
        13'd4357: m_out<=8'b11100010;
        13'd4358: m_out<=8'b00001100;
        13'd4359: m_out<=8'b00100001;
        13'd4360: m_out<=8'b11110101;
        13'd4361: m_out<=8'b00000110;
        13'd4362: m_out<=8'b00111001;
        13'd4363: m_out<=8'b11111011;
        13'd4364: m_out<=8'b00101011;
        13'd4365: m_out<=8'b00010001;
        13'd4366: m_out<=8'b11110001;
        13'd4367: m_out<=8'b11111111;
        13'd4368: m_out<=8'b00011101;
        13'd4369: m_out<=8'b00100001;
        13'd4370: m_out<=8'b11100110;
        13'd4371: m_out<=8'b11011101;
        13'd4372: m_out<=8'b11100000;
        13'd4373: m_out<=8'b11001010;
        13'd4374: m_out<=8'b00000000;
        13'd4375: m_out<=8'b00010100;
        13'd4376: m_out<=8'b00011111;
        13'd4377: m_out<=8'b11110001;
        13'd4378: m_out<=8'b11101000;
        13'd4379: m_out<=8'b00001000;
        13'd4380: m_out<=8'b00000001;
        13'd4381: m_out<=8'b00010110;
        13'd4382: m_out<=8'b00001011;
        13'd4383: m_out<=8'b00100010;
        13'd4384: m_out<=8'b00001110;
        13'd4385: m_out<=8'b11110111;
        13'd4386: m_out<=8'b11110111;
        13'd4387: m_out<=8'b11101010;
        13'd4388: m_out<=8'b00011101;
        13'd4389: m_out<=8'b00011000;
        13'd4390: m_out<=8'b00001000;
        13'd4391: m_out<=8'b11110001;
        13'd4392: m_out<=8'b11000000;
        13'd4393: m_out<=8'b11111111;
        13'd4394: m_out<=8'b00011101;
        13'd4395: m_out<=8'b00011110;
        13'd4396: m_out<=8'b00011000;
        13'd4397: m_out<=8'b11100110;
        13'd4398: m_out<=8'b00010011;
        13'd4399: m_out<=8'b00011101;
        13'd4400: m_out<=8'b11110111;
        13'd4401: m_out<=8'b11110110;
        13'd4402: m_out<=8'b11101010;
        13'd4403: m_out<=8'b11111101;
        13'd4404: m_out<=8'b11111110;
        13'd4405: m_out<=8'b00001110;
        13'd4406: m_out<=8'b00000111;
        13'd4407: m_out<=8'b11100111;
        13'd4408: m_out<=8'b11010100;
        13'd4409: m_out<=8'b11011101;
        13'd4410: m_out<=8'b11100100;
        13'd4411: m_out<=8'b00010111;
        13'd4412: m_out<=8'b11100011;
        13'd4413: m_out<=8'b00001001;
        13'd4414: m_out<=8'b00001010;
        13'd4415: m_out<=8'b11100110;
        13'd4416: m_out<=8'b00000010;
        13'd4417: m_out<=8'b00001011;
        13'd4418: m_out<=8'b11111101;
        13'd4419: m_out<=8'b11111011;
        13'd4420: m_out<=8'b11111101;
        13'd4421: m_out<=8'b00001111;
        13'd4422: m_out<=8'b00100000;
        13'd4423: m_out<=8'b00011000;
        13'd4424: m_out<=8'b00110001;
        13'd4425: m_out<=8'b11100100;
        13'd4426: m_out<=8'b00000110;
        13'd4427: m_out<=8'b11101111;
        13'd4428: m_out<=8'b10111101;
        13'd4429: m_out<=8'b00001011;
        13'd4430: m_out<=8'b00001100;
        13'd4431: m_out<=8'b11110011;
        13'd4432: m_out<=8'b11101001;
        13'd4433: m_out<=8'b11100100;
        13'd4434: m_out<=8'b00100010;
        13'd4435: m_out<=8'b00001000;
        13'd4436: m_out<=8'b00001011;
        13'd4437: m_out<=8'b00001101;
        13'd4438: m_out<=8'b11111110;
        13'd4439: m_out<=8'b11101111;
        13'd4440: m_out<=8'b11110000;
        13'd4441: m_out<=8'b11111000;
        13'd4442: m_out<=8'b11010111;
        13'd4443: m_out<=8'b00010110;
        13'd4444: m_out<=8'b00111110;
        13'd4445: m_out<=8'b00001101;
        13'd4446: m_out<=8'b00000101;
        13'd4447: m_out<=8'b00000111;
        13'd4448: m_out<=8'b11110000;
        13'd4449: m_out<=8'b11110101;
        13'd4450: m_out<=8'b00001011;
        13'd4451: m_out<=8'b11100010;
        13'd4452: m_out<=8'b11110101;
        13'd4453: m_out<=8'b11100100;
        13'd4454: m_out<=8'b00101001;
        13'd4455: m_out<=8'b00001111;
        13'd4456: m_out<=8'b11101101;
        13'd4457: m_out<=8'b00001101;
        13'd4458: m_out<=8'b00000110;
        13'd4459: m_out<=8'b11100000;
        13'd4460: m_out<=8'b11110100;
        13'd4461: m_out<=8'b00001100;
        13'd4462: m_out<=8'b11100001;
        13'd4463: m_out<=8'b11111101;
        13'd4464: m_out<=8'b11011010;
        13'd4465: m_out<=8'b00010011;
        13'd4466: m_out<=8'b00000100;
        13'd4467: m_out<=8'b11011001;
        13'd4468: m_out<=8'b11110110;
        13'd4469: m_out<=8'b11110100;
        13'd4470: m_out<=8'b00001111;
        13'd4471: m_out<=8'b00001110;
        13'd4472: m_out<=8'b11111101;
        13'd4473: m_out<=8'b00001001;
        13'd4474: m_out<=8'b11101101;
        13'd4475: m_out<=8'b11110100;
        13'd4476: m_out<=8'b00010010;
        13'd4477: m_out<=8'b00010010;
        13'd4478: m_out<=8'b00101101;
        13'd4479: m_out<=8'b11101111;
        13'd4480: m_out<=8'b00000100;
        13'd4481: m_out<=8'b11110001;
        13'd4482: m_out<=8'b11010101;
        13'd4483: m_out<=8'b11101000;
        13'd4484: m_out<=8'b11011100;
        13'd4485: m_out<=8'b11101101;
        13'd4486: m_out<=8'b00110011;
        13'd4487: m_out<=8'b00011101;
        13'd4488: m_out<=8'b00001001;
        13'd4489: m_out<=8'b00001101;
        13'd4490: m_out<=8'b11010110;
        13'd4491: m_out<=8'b00010001;
        13'd4492: m_out<=8'b11101000;
        13'd4493: m_out<=8'b00101000;
        13'd4494: m_out<=8'b00010100;
        13'd4495: m_out<=8'b11111001;
        13'd4496: m_out<=8'b00101010;
        13'd4497: m_out<=8'b00001100;
        13'd4498: m_out<=8'b00011011;
        13'd4499: m_out<=8'b00000000;
        13'd4500: m_out<=8'b11100001;
        13'd4501: m_out<=8'b11101011;
        13'd4502: m_out<=8'b11110011;
        13'd4503: m_out<=8'b00001010;
        13'd4504: m_out<=8'b11001011;
        13'd4505: m_out<=8'b11111111;
        13'd4506: m_out<=8'b00100111;
        13'd4507: m_out<=8'b00001000;
        13'd4508: m_out<=8'b11110111;
        13'd4509: m_out<=8'b00001110;
        13'd4510: m_out<=8'b11111100;
        13'd4511: m_out<=8'b11100101;
        13'd4512: m_out<=8'b00000001;
        13'd4513: m_out<=8'b00000000;
        13'd4514: m_out<=8'b00010001;
        13'd4515: m_out<=8'b11111010;
        13'd4516: m_out<=8'b11101111;
        13'd4517: m_out<=8'b11100011;
        13'd4518: m_out<=8'b11101110;
        13'd4519: m_out<=8'b00011100;
        13'd4520: m_out<=8'b00100100;
        13'd4521: m_out<=8'b00011100;
        13'd4522: m_out<=8'b11000101;
        13'd4523: m_out<=8'b11111100;
        13'd4524: m_out<=8'b00001100;
        13'd4525: m_out<=8'b11111001;
        13'd4526: m_out<=8'b11100111;
        13'd4527: m_out<=8'b11011000;
        13'd4528: m_out<=8'b00001111;
        13'd4529: m_out<=8'b00000000;
        13'd4530: m_out<=8'b11111001;
        13'd4531: m_out<=8'b11101111;
        13'd4532: m_out<=8'b00101101;
        13'd4533: m_out<=8'b11100111;
        13'd4534: m_out<=8'b00011110;
        13'd4535: m_out<=8'b11111010;
        13'd4536: m_out<=8'b11101100;
        13'd4537: m_out<=8'b00100110;
        13'd4538: m_out<=8'b00000100;
        13'd4539: m_out<=8'b11111111;
        13'd4540: m_out<=8'b11001111;
        13'd4541: m_out<=8'b00001011;
        13'd4542: m_out<=8'b00000001;
        13'd4543: m_out<=8'b11110010;
        13'd4544: m_out<=8'b11101000;
        13'd4545: m_out<=8'b00010010;
        13'd4546: m_out<=8'b00010011;
        13'd4547: m_out<=8'b11100011;
        13'd4548: m_out<=8'b00010000;
        13'd4549: m_out<=8'b00000000;
        13'd4550: m_out<=8'b11110101;
        13'd4551: m_out<=8'b00010101;
        13'd4552: m_out<=8'b11110100;
        13'd4553: m_out<=8'b00001011;
        13'd4554: m_out<=8'b11110100;
        13'd4555: m_out<=8'b11111010;
        13'd4556: m_out<=8'b11100011;
        13'd4557: m_out<=8'b00001001;
        13'd4558: m_out<=8'b00000111;
        13'd4559: m_out<=8'b00000110;
        13'd4560: m_out<=8'b11111010;
        13'd4561: m_out<=8'b11111010;
        13'd4562: m_out<=8'b11101101;
        13'd4563: m_out<=8'b00100100;
        13'd4564: m_out<=8'b00000010;
        13'd4565: m_out<=8'b00001101;
        13'd4566: m_out<=8'b11101110;
        13'd4567: m_out<=8'b00011010;
        13'd4568: m_out<=8'b11011011;
        13'd4569: m_out<=8'b00001010;
        13'd4570: m_out<=8'b00000100;
        13'd4571: m_out<=8'b00101100;
        13'd4572: m_out<=8'b11111100;
        13'd4573: m_out<=8'b11110000;
        13'd4574: m_out<=8'b11000110;
        13'd4575: m_out<=8'b11011011;
        13'd4576: m_out<=8'b01000100;
        13'd4577: m_out<=8'b11010011;
        13'd4578: m_out<=8'b11100111;
        13'd4579: m_out<=8'b00010110;
        13'd4580: m_out<=8'b11110011;
        13'd4581: m_out<=8'b11100100;
        13'd4582: m_out<=8'b00010110;
        13'd4583: m_out<=8'b11110000;
        13'd4584: m_out<=8'b11010010;
        13'd4585: m_out<=8'b11101011;
        13'd4586: m_out<=8'b11111010;
        13'd4587: m_out<=8'b11010011;
        13'd4588: m_out<=8'b00011100;
        13'd4589: m_out<=8'b00000000;
        13'd4590: m_out<=8'b11110001;
        13'd4591: m_out<=8'b11101011;
        13'd4592: m_out<=8'b11111011;
        13'd4593: m_out<=8'b00011101;
        13'd4594: m_out<=8'b11100001;
        13'd4595: m_out<=8'b00010011;
        13'd4596: m_out<=8'b00001110;
        13'd4597: m_out<=8'b11100010;
        13'd4598: m_out<=8'b11111101;
        13'd4599: m_out<=8'b11100001;
        13'd4600: m_out<=8'b00001110;
        13'd4601: m_out<=8'b00001000;
        13'd4602: m_out<=8'b11111111;
        13'd4603: m_out<=8'b11000010;
        13'd4604: m_out<=8'b00001001;
        13'd4605: m_out<=8'b00000111;
        13'd4606: m_out<=8'b00001001;
        13'd4607: m_out<=8'b00001111;
        13'd4608: m_out<=8'b11111011;
        13'd4609: m_out<=8'b11110101;
        13'd4610: m_out<=8'b11110001;
        13'd4611: m_out<=8'b11101010;
        13'd4612: m_out<=8'b11101101;
        13'd4613: m_out<=8'b11011110;
        13'd4614: m_out<=8'b11000110;
        13'd4615: m_out<=8'b00001110;
        13'd4616: m_out<=8'b11001011;
        13'd4617: m_out<=8'b00000100;
        13'd4618: m_out<=8'b11101100;
        13'd4619: m_out<=8'b11111100;
        13'd4620: m_out<=8'b00111000;
        13'd4621: m_out<=8'b00000001;
        13'd4622: m_out<=8'b00000101;
        13'd4623: m_out<=8'b00000000;
        13'd4624: m_out<=8'b00100110;
        13'd4625: m_out<=8'b11010110;
        13'd4626: m_out<=8'b01001011;
        13'd4627: m_out<=8'b00110000;
        13'd4628: m_out<=8'b11101101;
        13'd4629: m_out<=8'b00010110;
        13'd4630: m_out<=8'b11111111;
        13'd4631: m_out<=8'b11101110;
        13'd4632: m_out<=8'b11111111;
        13'd4633: m_out<=8'b00010101;
        13'd4634: m_out<=8'b00011101;
        13'd4635: m_out<=8'b00000110;
        13'd4636: m_out<=8'b00010100;
        13'd4637: m_out<=8'b00001111;
        13'd4638: m_out<=8'b11101011;
        13'd4639: m_out<=8'b11110111;
        13'd4640: m_out<=8'b11101001;
        13'd4641: m_out<=8'b11111010;
        13'd4642: m_out<=8'b00001110;
        13'd4643: m_out<=8'b00101000;
        13'd4644: m_out<=8'b00101111;
        13'd4645: m_out<=8'b00010111;
        13'd4646: m_out<=8'b11101000;
        13'd4647: m_out<=8'b11111000;
        13'd4648: m_out<=8'b11110010;
        13'd4649: m_out<=8'b11111001;
        13'd4650: m_out<=8'b00010010;
        13'd4651: m_out<=8'b11101101;
        13'd4652: m_out<=8'b00010000;
        13'd4653: m_out<=8'b00011101;
        13'd4654: m_out<=8'b00000011;
        13'd4655: m_out<=8'b11111110;
        13'd4656: m_out<=8'b11111010;
        13'd4657: m_out<=8'b11101010;
        13'd4658: m_out<=8'b11101111;
        13'd4659: m_out<=8'b11110100;
        13'd4660: m_out<=8'b11101101;
        13'd4661: m_out<=8'b00110001;
        13'd4662: m_out<=8'b11011111;
        13'd4663: m_out<=8'b11001101;
        13'd4664: m_out<=8'b11100100;
        13'd4665: m_out<=8'b11110011;
        13'd4666: m_out<=8'b00001101;
        13'd4667: m_out<=8'b00000011;
        13'd4668: m_out<=8'b11110110;
        13'd4669: m_out<=8'b00101011;
        13'd4670: m_out<=8'b00001011;
        13'd4671: m_out<=8'b11011111;
        13'd4672: m_out<=8'b11111100;
        13'd4673: m_out<=8'b00101000;
        13'd4674: m_out<=8'b00000101;
        13'd4675: m_out<=8'b11100100;
        13'd4676: m_out<=8'b00000011;
        13'd4677: m_out<=8'b11110001;
        13'd4678: m_out<=8'b11110000;
        13'd4679: m_out<=8'b00000100;
        13'd4680: m_out<=8'b11110000;
        13'd4681: m_out<=8'b00110011;
        13'd4682: m_out<=8'b00011100;
        13'd4683: m_out<=8'b00001101;
        13'd4684: m_out<=8'b00011011;
        13'd4685: m_out<=8'b11111101;
        13'd4686: m_out<=8'b00011000;
        13'd4687: m_out<=8'b00001001;
        13'd4688: m_out<=8'b00001101;
        13'd4689: m_out<=8'b11001000;
        13'd4690: m_out<=8'b00001010;
        13'd4691: m_out<=8'b00000011;
        13'd4692: m_out<=8'b00100001;
        13'd4693: m_out<=8'b00000111;
        13'd4694: m_out<=8'b00000001;
        13'd4695: m_out<=8'b00000000;
        13'd4696: m_out<=8'b00000111;
        13'd4697: m_out<=8'b11101010;
        13'd4698: m_out<=8'b11110000;
        13'd4699: m_out<=8'b11101101;
        13'd4700: m_out<=8'b00010011;
        13'd4701: m_out<=8'b00000011;
        13'd4702: m_out<=8'b11101001;
        13'd4703: m_out<=8'b11101111;
        13'd4704: m_out<=8'b11100110;
        13'd4705: m_out<=8'b00010100;
        13'd4706: m_out<=8'b11101111;
        13'd4707: m_out<=8'b00000010;
        13'd4708: m_out<=8'b00010001;
        13'd4709: m_out<=8'b11110111;
        13'd4710: m_out<=8'b11100111;
        13'd4711: m_out<=8'b11111011;
        13'd4712: m_out<=8'b00100101;
        13'd4713: m_out<=8'b00011110;
        13'd4714: m_out<=8'b00001100;
        13'd4715: m_out<=8'b00010110;
        13'd4716: m_out<=8'b00101100;
        13'd4717: m_out<=8'b00010011;
        13'd4718: m_out<=8'b00000000;
        13'd4719: m_out<=8'b00001100;
        13'd4720: m_out<=8'b11010100;
        13'd4721: m_out<=8'b11100111;
        13'd4722: m_out<=8'b11001110;
        13'd4723: m_out<=8'b00001100;
        13'd4724: m_out<=8'b00110001;
        13'd4725: m_out<=8'b11110011;
        13'd4726: m_out<=8'b00100101;
        13'd4727: m_out<=8'b00001001;
        13'd4728: m_out<=8'b00010101;
        13'd4729: m_out<=8'b00010000;
        13'd4730: m_out<=8'b11011111;
        13'd4731: m_out<=8'b11011010;
        13'd4732: m_out<=8'b00000110;
        13'd4733: m_out<=8'b11010101;
        13'd4734: m_out<=8'b00010100;
        13'd4735: m_out<=8'b00001001;
        13'd4736: m_out<=8'b11101000;
        13'd4737: m_out<=8'b00100001;
        13'd4738: m_out<=8'b11101111;
        13'd4739: m_out<=8'b00110111;
        13'd4740: m_out<=8'b00010110;
        13'd4741: m_out<=8'b11010000;
        13'd4742: m_out<=8'b11011111;
        13'd4743: m_out<=8'b11111000;
        13'd4744: m_out<=8'b11111101;
        13'd4745: m_out<=8'b00001100;
        13'd4746: m_out<=8'b00000100;
        13'd4747: m_out<=8'b11001010;
        13'd4748: m_out<=8'b11111010;
        13'd4749: m_out<=8'b00010101;
        13'd4750: m_out<=8'b00010010;
        13'd4751: m_out<=8'b00010100;
        13'd4752: m_out<=8'b00111000;
        13'd4753: m_out<=8'b00010101;
        13'd4754: m_out<=8'b11111001;
        13'd4755: m_out<=8'b00110100;
        13'd4756: m_out<=8'b11111110;
        13'd4757: m_out<=8'b11111110;
        13'd4758: m_out<=8'b11110111;
        13'd4759: m_out<=8'b11110011;
        13'd4760: m_out<=8'b11111101;
        13'd4761: m_out<=8'b11101110;
        13'd4762: m_out<=8'b11011111;
        13'd4763: m_out<=8'b00001100;
        13'd4764: m_out<=8'b00100000;
        13'd4765: m_out<=8'b00011011;
        13'd4766: m_out<=8'b00010110;
        13'd4767: m_out<=8'b11000100;
        13'd4768: m_out<=8'b11101011;
        13'd4769: m_out<=8'b00111100;
        13'd4770: m_out<=8'b11011100;
        13'd4771: m_out<=8'b00011011;
        13'd4772: m_out<=8'b11101101;
        13'd4773: m_out<=8'b11111000;
        13'd4774: m_out<=8'b11110110;
        13'd4775: m_out<=8'b00110110;
        13'd4776: m_out<=8'b00000100;
        13'd4777: m_out<=8'b00001111;
        13'd4778: m_out<=8'b00010010;
        13'd4779: m_out<=8'b00100001;
        13'd4780: m_out<=8'b00010110;
        13'd4781: m_out<=8'b00010000;
        13'd4782: m_out<=8'b00001100;
        13'd4783: m_out<=8'b11111110;
        13'd4784: m_out<=8'b11111101;
        13'd4785: m_out<=8'b00100000;
        13'd4786: m_out<=8'b11000110;
        13'd4787: m_out<=8'b00100010;
        13'd4788: m_out<=8'b00011101;
        13'd4789: m_out<=8'b00000001;
        13'd4790: m_out<=8'b00111110;
        13'd4791: m_out<=8'b11111011;
        13'd4792: m_out<=8'b11111010;
        13'd4793: m_out<=8'b11101100;
        13'd4794: m_out<=8'b00011111;
        13'd4795: m_out<=8'b00000001;
        13'd4796: m_out<=8'b00000011;
        13'd4797: m_out<=8'b00000100;
        13'd4798: m_out<=8'b11111010;
        13'd4799: m_out<=8'b11101101;
        13'd4800: m_out<=8'b00000010;
        13'd4801: m_out<=8'b00011001;
        13'd4802: m_out<=8'b00000010;
        13'd4803: m_out<=8'b11010001;
        13'd4804: m_out<=8'b11111101;
        13'd4805: m_out<=8'b11100001;
        13'd4806: m_out<=8'b11111011;
        13'd4807: m_out<=8'b11110000;
        13'd4808: m_out<=8'b11100010;
        13'd4809: m_out<=8'b11110111;
        13'd4810: m_out<=8'b00011110;
        13'd4811: m_out<=8'b00010001;
        13'd4812: m_out<=8'b00001010;
        13'd4813: m_out<=8'b00000111;
        13'd4814: m_out<=8'b00101000;
        13'd4815: m_out<=8'b00111111;
        13'd4816: m_out<=8'b11101100;
        13'd4817: m_out<=8'b11001100;
        13'd4818: m_out<=8'b11111011;
        13'd4819: m_out<=8'b00001001;
        13'd4820: m_out<=8'b11101011;
        13'd4821: m_out<=8'b00011101;
        13'd4822: m_out<=8'b00010111;
        13'd4823: m_out<=8'b11101101;
        13'd4824: m_out<=8'b00000000;
        13'd4825: m_out<=8'b00011110;
        13'd4826: m_out<=8'b11110001;
        13'd4827: m_out<=8'b11101011;
        13'd4828: m_out<=8'b11111000;
        13'd4829: m_out<=8'b00110001;
        13'd4830: m_out<=8'b11011111;
        13'd4831: m_out<=8'b11111000;
        13'd4832: m_out<=8'b11111100;
        13'd4833: m_out<=8'b00001000;
        13'd4834: m_out<=8'b00001100;
        13'd4835: m_out<=8'b00101000;
        13'd4836: m_out<=8'b11111111;
        13'd4837: m_out<=8'b11110110;
        13'd4838: m_out<=8'b00001111;
        13'd4839: m_out<=8'b00100011;
        13'd4840: m_out<=8'b11110001;
        13'd4841: m_out<=8'b00010001;
        13'd4842: m_out<=8'b00000101;
        13'd4843: m_out<=8'b11110111;
        13'd4844: m_out<=8'b11110111;
        13'd4845: m_out<=8'b00010100;
        13'd4846: m_out<=8'b00100000;
        13'd4847: m_out<=8'b01000001;
        13'd4848: m_out<=8'b00010000;
        13'd4849: m_out<=8'b00010100;
        13'd4850: m_out<=8'b11110001;
        13'd4851: m_out<=8'b11110001;
        13'd4852: m_out<=8'b11100111;
        13'd4853: m_out<=8'b11111111;
        13'd4854: m_out<=8'b00100111;
        13'd4855: m_out<=8'b11110100;
        13'd4856: m_out<=8'b11111010;
        13'd4857: m_out<=8'b00000010;
        13'd4858: m_out<=8'b00000000;
        13'd4859: m_out<=8'b11111110;
        13'd4860: m_out<=8'b01000111;
        13'd4861: m_out<=8'b11101111;
        13'd4862: m_out<=8'b00000110;
        13'd4863: m_out<=8'b00000011;
        13'd4864: m_out<=8'b11111010;
        13'd4865: m_out<=8'b11110000;
        13'd4866: m_out<=8'b00110000;
        13'd4867: m_out<=8'b11111100;
        13'd4868: m_out<=8'b00101010;
        13'd4869: m_out<=8'b00001111;
        13'd4870: m_out<=8'b00000000;
        13'd4871: m_out<=8'b00110011;
        13'd4872: m_out<=8'b11111111;
        13'd4873: m_out<=8'b11100001;
        13'd4874: m_out<=8'b00000100;
        13'd4875: m_out<=8'b00010101;
        13'd4876: m_out<=8'b11100111;
        13'd4877: m_out<=8'b11110110;
        13'd4878: m_out<=8'b11111010;
        13'd4879: m_out<=8'b11101110;
        13'd4880: m_out<=8'b11110111;
        13'd4881: m_out<=8'b11110110;
        13'd4882: m_out<=8'b00010010;
        13'd4883: m_out<=8'b00110111;
        13'd4884: m_out<=8'b11010111;
        13'd4885: m_out<=8'b11010111;
        13'd4886: m_out<=8'b00011101;
        13'd4887: m_out<=8'b11011001;
        13'd4888: m_out<=8'b11111111;
        13'd4889: m_out<=8'b00001100;
        13'd4890: m_out<=8'b11110010;
        13'd4891: m_out<=8'b11101110;
        13'd4892: m_out<=8'b00001001;
        13'd4893: m_out<=8'b11110100;
        13'd4894: m_out<=8'b00010101;
        13'd4895: m_out<=8'b11110111;
        13'd4896: m_out<=8'b11111111;
        13'd4897: m_out<=8'b00110010;
        13'd4898: m_out<=8'b11000100;
        13'd4899: m_out<=8'b00000010;
        13'd4900: m_out<=8'b11011110;
        13'd4901: m_out<=8'b00010010;
        13'd4902: m_out<=8'b00010011;
        13'd4903: m_out<=8'b11100010;
        13'd4904: m_out<=8'b11101001;
        13'd4905: m_out<=8'b00010110;
        13'd4906: m_out<=8'b11101111;
        13'd4907: m_out<=8'b00011100;
        13'd4908: m_out<=8'b11011101;
        13'd4909: m_out<=8'b11110010;
        13'd4910: m_out<=8'b11101011;
        13'd4911: m_out<=8'b00101001;
        13'd4912: m_out<=8'b00001010;
        13'd4913: m_out<=8'b00010000;
        13'd4914: m_out<=8'b00000011;
        13'd4915: m_out<=8'b00000110;
        13'd4916: m_out<=8'b00000000;
        13'd4917: m_out<=8'b00000110;
        13'd4918: m_out<=8'b11101100;
        13'd4919: m_out<=8'b00000000;
        13'd4920: m_out<=8'b00011001;
        13'd4921: m_out<=8'b11110011;
        13'd4922: m_out<=8'b11101001;
        13'd4923: m_out<=8'b11101110;
        13'd4924: m_out<=8'b00001110;
        13'd4925: m_out<=8'b11111100;
        13'd4926: m_out<=8'b00010110;
        13'd4927: m_out<=8'b00011010;
        13'd4928: m_out<=8'b00010101;
        13'd4929: m_out<=8'b11100011;
        13'd4930: m_out<=8'b11011111;
        13'd4931: m_out<=8'b00010100;
        13'd4932: m_out<=8'b11111000;
        13'd4933: m_out<=8'b11111110;
        13'd4934: m_out<=8'b11110001;
        13'd4935: m_out<=8'b00010010;
        13'd4936: m_out<=8'b11101111;
        13'd4937: m_out<=8'b11101001;
        13'd4938: m_out<=8'b11111100;
        13'd4939: m_out<=8'b11110110;
        13'd4940: m_out<=8'b00101011;
        13'd4941: m_out<=8'b00001011;
        13'd4942: m_out<=8'b00011101;
        13'd4943: m_out<=8'b11100111;
        13'd4944: m_out<=8'b00010000;
        13'd4945: m_out<=8'b11110101;
        13'd4946: m_out<=8'b00010010;
        13'd4947: m_out<=8'b11110000;
        13'd4948: m_out<=8'b11101100;
        13'd4949: m_out<=8'b11001110;
        13'd4950: m_out<=8'b00000011;
        13'd4951: m_out<=8'b11110111;
        13'd4952: m_out<=8'b11111001;
        13'd4953: m_out<=8'b11010110;
        13'd4954: m_out<=8'b11111010;
        13'd4955: m_out<=8'b00110100;
        13'd4956: m_out<=8'b11101001;
        13'd4957: m_out<=8'b11111001;
        13'd4958: m_out<=8'b00100001;
        13'd4959: m_out<=8'b00111001;
        13'd4960: m_out<=8'b11010110;
        13'd4961: m_out<=8'b11100010;
        13'd4962: m_out<=8'b11111100;
        13'd4963: m_out<=8'b11110110;
        13'd4964: m_out<=8'b11100000;
        13'd4965: m_out<=8'b00010110;
        13'd4966: m_out<=8'b11110110;
        13'd4967: m_out<=8'b00011110;
        13'd4968: m_out<=8'b11011100;
        13'd4969: m_out<=8'b00000010;
        13'd4970: m_out<=8'b11010000;
        13'd4971: m_out<=8'b00010000;
        13'd4972: m_out<=8'b00100000;
        13'd4973: m_out<=8'b00000001;
        13'd4974: m_out<=8'b00110010;
        13'd4975: m_out<=8'b00110111;
        13'd4976: m_out<=8'b11100010;
        13'd4977: m_out<=8'b00101011;
        13'd4978: m_out<=8'b00011001;
        13'd4979: m_out<=8'b00000100;
        13'd4980: m_out<=8'b11111000;
        13'd4981: m_out<=8'b11000111;
        13'd4982: m_out<=8'b11100010;
        13'd4983: m_out<=8'b11111110;
        13'd4984: m_out<=8'b00000101;
        13'd4985: m_out<=8'b11100101;
        13'd4986: m_out<=8'b00010011;
        13'd4987: m_out<=8'b11101101;
        13'd4988: m_out<=8'b00010010;
        13'd4989: m_out<=8'b00010011;
        13'd4990: m_out<=8'b11111001;
        13'd4991: m_out<=8'b11111100;
        13'd4992: m_out<=8'b10111011;
        13'd4993: m_out<=8'b11110010;
        13'd4994: m_out<=8'b00010000;
        13'd4995: m_out<=8'b11110111;
        13'd4996: m_out<=8'b11110100;
        13'd4997: m_out<=8'b00010000;
        13'd4998: m_out<=8'b11100100;
        13'd4999: m_out<=8'b11100111;
        default: m_out <=8'b0;
    endcase
assign out = m_out;
endmodule
