module IOTProject(
	input clk
);

	mySystem u0 (
		.clk_clk (clk)  // clk.clk
	);



endmodule
