module generator(
	output[7:0] rec,

	output rst,
	output ena,
	output clk
);

reg[7:0] sig;
reg m_rst;
reg m_ena;
reg m_clk;


always@(*) begin
	m_clk = 0;
	#500;
	m_clk = ~clk;
	#1000;
	m_clk = ~clk;
end

initial begin
	sig = 8'b11100100;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b01000110;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00111000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b11001000;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b10111111;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11000010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00111000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b01100001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b10111101;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b10111110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00111011;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00111001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b10111111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00111011;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b01001001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b01000011;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b01000111;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11000010;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b10110010;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00111000;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b01001010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00111101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b10111011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00111101;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b10111101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b01001100;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00111111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b10110110;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b01001011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b01001001;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00111100;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b01010101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b01000001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b10110001;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b01000010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b10110001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11000001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00111000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b10111111;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b00111000;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00111011;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00110010;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b10111011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00111010;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11000011;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b10111011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b10111010;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b10111010;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b00111111;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00110010;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b00111001;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11001001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b01000001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b11001001;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b00111101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00111010;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b10101100;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00110010;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11001001;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00111001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11000010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b01000001;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b01000100;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b10111111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b01000100;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11001000;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b01000100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00110010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00111000;
#1000;
sig = 8'b00111011;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b01000000;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11000011;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00110010;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00111001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b10111100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11001001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11000000;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b10111101;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00111010;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b01000111;
#1000;
sig = 8'b01010100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b01000011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b10011111;
#1000;
sig = 8'b10011111;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b10111101;
#1000;
sig = 8'b10100010;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00111010;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b10111100;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00110010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11000011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b01000000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b01000110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b01000011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00111101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b01000101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11001000;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b01011011;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b10111100;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00111011;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b01000010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11001001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b10111100;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b01001000;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00101110;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b01011010;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00111100;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b10101110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00111011;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b10111101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b11000001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00111101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11000011;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b00111010;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00110101;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11001001;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00111111;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00111001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b10101101;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b01001001;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00111001;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11000000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b10111101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11000101;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11011000;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00101101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11001111;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00100100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b11011011;
#1000;
sig = 8'b01000100;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11010010;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11010011;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11000010;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11001011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00111000;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00100110;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b01001011;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00101111;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11001101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00011000;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00001101;
#1000;
sig = 8'b11001000;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b11101010;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11100110;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00101100;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11010100;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b00100101;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11011010;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11010101;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101000;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11001010;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00111000;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00111100;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00011011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00110110;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b11000110;
#1000;
sig = 8'b00100010;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00111110;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00011111;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11010001;
#1000;
sig = 8'b11111101;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00000111;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b00111111;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11001100;
#1000;
sig = 8'b11111011;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b00010111;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b00110001;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00001000;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b00101000;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00100011;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00010001;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b01000001;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00100111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b01000111;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b00110000;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00101010;
#1000;
sig = 8'b00001111;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00110011;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b11100001;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b11010111;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11011001;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00001100;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00001001;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111111;
#1000;
sig = 8'b00110010;
#1000;
sig = 8'b11000100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11011110;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b00011100;
#1000;
sig = 8'b11011101;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b11101011;
#1000;
sig = 8'b00101001;
#1000;
sig = 8'b00001010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00000110;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b00000000;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b11110011;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11101110;
#1000;
sig = 8'b00001110;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b00011010;
#1000;
sig = 8'b00010101;
#1000;
sig = 8'b11100011;
#1000;
sig = 8'b11011111;
#1000;
sig = 8'b00010100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b11110001;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11101111;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b00001011;
#1000;
sig = 8'b00011101;
#1000;
sig = 8'b11100111;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11110101;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b11110000;
#1000;
sig = 8'b11101100;
#1000;
sig = 8'b11001110;
#1000;
sig = 8'b00000011;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b11111010;
#1000;
sig = 8'b00110100;
#1000;
sig = 8'b11101001;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b00100001;
#1000;
sig = 8'b00111001;
#1000;
sig = 8'b11010110;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b11100000;
#1000;
sig = 8'b00010110;
#1000;
sig = 8'b11110110;
#1000;
sig = 8'b00011110;
#1000;
sig = 8'b11011100;
#1000;
sig = 8'b00000010;
#1000;
sig = 8'b11010000;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b00100000;
#1000;
sig = 8'b00000001;
#1000;
sig = 8'b00110010;
#1000;
sig = 8'b00110111;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b00101011;
#1000;
sig = 8'b00011001;
#1000;
sig = 8'b00000100;
#1000;
sig = 8'b11111000;
#1000;
sig = 8'b11000111;
#1000;
sig = 8'b11100010;
#1000;
sig = 8'b11111110;
#1000;
sig = 8'b00000101;
#1000;
sig = 8'b11100101;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11101101;
#1000;
sig = 8'b00010010;
#1000;
sig = 8'b00010011;
#1000;
sig = 8'b11111001;
#1000;
sig = 8'b11111100;
#1000;
sig = 8'b10111011;
#1000;
sig = 8'b11110010;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11110111;
#1000;
sig = 8'b11110100;
#1000;
sig = 8'b00010000;
#1000;
sig = 8'b11100100;
#1000;
sig = 8'b11100111;
#1000;
$finish;
end

assign rec = sig;
assign rst = m_rst;
assign ena = m_ena;
assign clk = m_clk;

endmodule
