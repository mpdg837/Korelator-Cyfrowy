// mySystem.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module mySystem (
		input  wire       clk_clk,              //          clk.clk
		input  wire [3:0] inputin_keys,         //      inputin.keys
		output wire [3:0] inputin_leds,         //             .leds
		input  wire       reset_reset_n,        //        reset.reset_n
		output wire [3:0] sevensegment_output1, // sevensegment.output1
		output wire [7:0] sevensegment_output,  //             .output
		input  wire       uart_rx,              //         uart.rx
		output wire       uart_tx               //             .tx
	);

	wire  [31:0] cpu_data_master_readdata;                                   // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                                // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                                // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [14:0] cpu_data_master_address;                                    // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                 // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                       // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                      // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                  // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                            // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                         // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [14:0] cpu_instruction_master_address;                             // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                                // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         uart_fast_0_m1_waitrequest;                                 // mm_interconnect_0:UART_Fast_0_m1_waitrequest -> UART_Fast_0:avm_m1_waitrequest
	wire  [31:0] uart_fast_0_m1_readdata;                                    // mm_interconnect_0:UART_Fast_0_m1_readdata -> UART_Fast_0:avm_m1_readdata
	wire         uart_fast_0_m1_read;                                        // UART_Fast_0:avm_m1_read -> mm_interconnect_0:UART_Fast_0_m1_read
	wire  [15:0] uart_fast_0_m1_address;                                     // UART_Fast_0:avm_m1_address -> mm_interconnect_0:UART_Fast_0_m1_address
	wire         uart_fast_0_m1_readdatavalid;                               // mm_interconnect_0:UART_Fast_0_m1_readdatavalid -> UART_Fast_0:avm_m1_readdatavalid
	wire         uart_fast_0_m1_write;                                       // UART_Fast_0:avm_m1_write -> mm_interconnect_0:UART_Fast_0_m1_write
	wire  [31:0] uart_fast_0_m1_writedata;                                   // UART_Fast_0:avm_m1_writedata -> mm_interconnect_0:UART_Fast_0_m1_writedata
	wire         conclover_0_m1_waitrequest;                                 // mm_interconnect_0:Conclover_0_m1_waitrequest -> Conclover_0:avm_m1_waitrequest
	wire  [31:0] conclover_0_m1_readdata;                                    // mm_interconnect_0:Conclover_0_m1_readdata -> Conclover_0:avm_m1_readdata
	wire         conclover_0_m1_read;                                        // Conclover_0:avm_m1_read -> mm_interconnect_0:Conclover_0_m1_read
	wire  [15:0] conclover_0_m1_address;                                     // Conclover_0:avm_m1_address -> mm_interconnect_0:Conclover_0_m1_address
	wire         conclover_0_m1_readdatavalid;                               // mm_interconnect_0:Conclover_0_m1_readdatavalid -> Conclover_0:avm_m1_readdatavalid
	wire         conclover_0_m1_write;                                       // Conclover_0:avm_m1_write -> mm_interconnect_0:Conclover_0_m1_write
	wire  [31:0] conclover_0_m1_writedata;                                   // Conclover_0:avm_m1_writedata -> mm_interconnect_0:Conclover_0_m1_writedata
	wire         mm_interconnect_0_debug_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:Debug_UART_avalon_jtag_slave_chipselect -> Debug_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_uart_avalon_jtag_slave_readdata;    // Debug_UART:av_readdata -> mm_interconnect_0:Debug_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_uart_avalon_jtag_slave_waitrequest; // Debug_UART:av_waitrequest -> mm_interconnect_0:Debug_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_uart_avalon_jtag_slave_address;     // mm_interconnect_0:Debug_UART_avalon_jtag_slave_address -> Debug_UART:av_address
	wire         mm_interconnect_0_debug_uart_avalon_jtag_slave_read;        // mm_interconnect_0:Debug_UART_avalon_jtag_slave_read -> Debug_UART:av_read_n
	wire         mm_interconnect_0_debug_uart_avalon_jtag_slave_write;       // mm_interconnect_0:Debug_UART_avalon_jtag_slave_write -> Debug_UART:av_write_n
	wire  [31:0] mm_interconnect_0_debug_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:Debug_UART_avalon_jtag_slave_writedata -> Debug_UART:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;             // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;          // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;          // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;              // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                 // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;           // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;            // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_seven_segment_display_s0_readdata;        // Seven_Segment_Display:avs_s0_readdata -> mm_interconnect_0:Seven_Segment_Display_s0_readdata
	wire   [4:0] mm_interconnect_0_seven_segment_display_s0_address;         // mm_interconnect_0:Seven_Segment_Display_s0_address -> Seven_Segment_Display:avs_s0_address
	wire         mm_interconnect_0_seven_segment_display_s0_read;            // mm_interconnect_0:Seven_Segment_Display_s0_read -> Seven_Segment_Display:avs_s0_read
	wire         mm_interconnect_0_seven_segment_display_s0_write;           // mm_interconnect_0:Seven_Segment_Display_s0_write -> Seven_Segment_Display:avs_s0_write
	wire  [31:0] mm_interconnect_0_seven_segment_display_s0_writedata;       // mm_interconnect_0:Seven_Segment_Display_s0_writedata -> Seven_Segment_Display:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_system_timer_s0_readdata;                 // System_Timer:avs_s0_readdata -> mm_interconnect_0:System_Timer_s0_readdata
	wire   [1:0] mm_interconnect_0_system_timer_s0_address;                  // mm_interconnect_0:System_Timer_s0_address -> System_Timer:avs_s0_address
	wire         mm_interconnect_0_system_timer_s0_read;                     // mm_interconnect_0:System_Timer_s0_read -> System_Timer:avs_s0_read
	wire         mm_interconnect_0_system_timer_s0_write;                    // mm_interconnect_0:System_Timer_s0_write -> System_Timer:avs_s0_write
	wire  [31:0] mm_interconnect_0_system_timer_s0_writedata;                // mm_interconnect_0:System_Timer_s0_writedata -> System_Timer:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_input_s0_readdata;                        // Input:avs_s0_readdata -> mm_interconnect_0:Input_s0_readdata
	wire   [3:0] mm_interconnect_0_input_s0_address;                         // mm_interconnect_0:Input_s0_address -> Input:avs_s0_address
	wire         mm_interconnect_0_input_s0_read;                            // mm_interconnect_0:Input_s0_read -> Input:avs_s0_read
	wire         mm_interconnect_0_input_s0_write;                           // mm_interconnect_0:Input_s0_write -> Input:avs_s0_write
	wire  [31:0] mm_interconnect_0_input_s0_writedata;                       // mm_interconnect_0:Input_s0_writedata -> Input:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_uart_fast_0_s0_readdata;                  // UART_Fast_0:avs_s0_readdata -> mm_interconnect_0:UART_Fast_0_s0_readdata
	wire   [2:0] mm_interconnect_0_uart_fast_0_s0_address;                   // mm_interconnect_0:UART_Fast_0_s0_address -> UART_Fast_0:avs_s0_address
	wire         mm_interconnect_0_uart_fast_0_s0_read;                      // mm_interconnect_0:UART_Fast_0_s0_read -> UART_Fast_0:avs_s0_read
	wire         mm_interconnect_0_uart_fast_0_s0_write;                     // mm_interconnect_0:UART_Fast_0_s0_write -> UART_Fast_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_uart_fast_0_s0_writedata;                 // mm_interconnect_0:UART_Fast_0_s0_writedata -> UART_Fast_0:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_conclover_0_s0_readdata;                  // Conclover_0:avs_s0_readdata -> mm_interconnect_0:Conclover_0_s0_readdata
	wire   [4:0] mm_interconnect_0_conclover_0_s0_address;                   // mm_interconnect_0:Conclover_0_s0_address -> Conclover_0:avs_s0_address
	wire         mm_interconnect_0_conclover_0_s0_read;                      // mm_interconnect_0:Conclover_0_s0_read -> Conclover_0:avs_s0_read
	wire         mm_interconnect_0_conclover_0_s0_write;                     // mm_interconnect_0:Conclover_0_s0_write -> Conclover_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_conclover_0_s0_writedata;                 // mm_interconnect_0:Conclover_0_s0_writedata -> Conclover_0:avs_s0_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                        // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                          // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                           // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                        // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                             // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                         // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                             // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         irq_mapper_receiver0_irq;                                   // Debug_UART:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_irq_irq;                                                // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [CPU:reset_n, Conclover_0:rsi_reset_n, Debug_UART:rst_n, Input:rsi_reset_n, RAM:reset, Seven_Segment_Display:rsi_reset_n, System_Timer:rsi_reset_n, UART_Fast_0:rsi_reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                              // CPU:debug_reset_request -> rst_controller:reset_in1

	mySystem_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	conclover conclover_0 (
		.csi_clk              (clk_clk),                                    // clock.clk
		.rsi_reset_n          (~rst_controller_reset_out_reset),            // reset.reset_n
		.avs_s0_write         (mm_interconnect_0_conclover_0_s0_write),     //    s0.write
		.avs_s0_read          (mm_interconnect_0_conclover_0_s0_read),      //      .read
		.avs_s0_address       (mm_interconnect_0_conclover_0_s0_address),   //      .address
		.avs_s0_writedata     (mm_interconnect_0_conclover_0_s0_writedata), //      .writedata
		.avs_s0_readdata      (mm_interconnect_0_conclover_0_s0_readdata),  //      .readdata
		.avm_m1_write         (conclover_0_m1_write),                       //    m1.write
		.avm_m1_read          (conclover_0_m1_read),                        //      .read
		.avm_m1_waitrequest   (conclover_0_m1_waitrequest),                 //      .waitrequest
		.avm_m1_readdatavalid (conclover_0_m1_readdatavalid),               //      .readdatavalid
		.avm_m1_address       (conclover_0_m1_address),                     //      .address
		.avm_m1_writedata     (conclover_0_m1_writedata),                   //      .writedata
		.avm_m1_readdata      (conclover_0_m1_readdata)                     //      .readdata
	);

	mySystem_Debug_UART debug_uart (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                            //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                    //               irq.irq
	);

	keyInput input_inst (
		.csi_clk          (clk_clk),                              //           clock.clk
		.rsi_reset_n      (~rst_controller_reset_out_reset),      //           reset.reset_n
		.avs_s0_write     (mm_interconnect_0_input_s0_write),     //              s0.write
		.avs_s0_read      (mm_interconnect_0_input_s0_read),      //                .read
		.avs_s0_address   (mm_interconnect_0_input_s0_address),   //                .address
		.avs_s0_writedata (mm_interconnect_0_input_s0_writedata), //                .writedata
		.avs_s0_readdata  (mm_interconnect_0_input_s0_readdata),  //                .readdata
		.in_key           (inputin_keys),                         // external_output.keys
		.out_led          (inputin_leds)                          //                .leds
	);

	mySystem_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	segmentDisplay seven_segment_display (
		.csi_clk          (clk_clk),                                              //           clock.clk
		.rsi_reset_n      (~rst_controller_reset_out_reset),                      //           reset.reset_n
		.avs_s0_write     (mm_interconnect_0_seven_segment_display_s0_write),     //              s0.write
		.avs_s0_read      (mm_interconnect_0_seven_segment_display_s0_read),      //                .read
		.avs_s0_address   (mm_interconnect_0_seven_segment_display_s0_address),   //                .address
		.avs_s0_writedata (mm_interconnect_0_seven_segment_display_s0_writedata), //                .writedata
		.avs_s0_readdata  (mm_interconnect_0_seven_segment_display_s0_readdata),  //                .readdata
		.out_dig          (sevensegment_output1),                                 // external_output.output1
		.out_segment      (sevensegment_output)                                   //                .output
	);

	timerModule system_timer (
		.csi_clk          (clk_clk),                                     // clock.clk
		.rsi_reset_n      (~rst_controller_reset_out_reset),             // reset.reset_n
		.avs_s0_write     (mm_interconnect_0_system_timer_s0_write),     //    s0.write
		.avs_s0_read      (mm_interconnect_0_system_timer_s0_read),      //      .read
		.avs_s0_address   (mm_interconnect_0_system_timer_s0_address),   //      .address
		.avs_s0_writedata (mm_interconnect_0_system_timer_s0_writedata), //      .writedata
		.avs_s0_readdata  (mm_interconnect_0_system_timer_s0_readdata)   //      .readdata
	);

	UART_Fast uart_fast_0 (
		.csi_clk              (clk_clk),                                    //       clock.clk
		.rsi_reset_n          (~rst_controller_reset_out_reset),            //       reset.reset_n
		.avs_s0_write         (mm_interconnect_0_uart_fast_0_s0_write),     //          s0.write
		.avs_s0_read          (mm_interconnect_0_uart_fast_0_s0_read),      //            .read
		.avs_s0_address       (mm_interconnect_0_uart_fast_0_s0_address),   //            .address
		.avs_s0_writedata     (mm_interconnect_0_uart_fast_0_s0_writedata), //            .writedata
		.avs_s0_readdata      (mm_interconnect_0_uart_fast_0_s0_readdata),  //            .readdata
		.avm_m1_write         (uart_fast_0_m1_write),                       //          m1.write
		.avm_m1_read          (uart_fast_0_m1_read),                        //            .read
		.avm_m1_waitrequest   (uart_fast_0_m1_waitrequest),                 //            .waitrequest
		.avm_m1_readdatavalid (uart_fast_0_m1_readdatavalid),               //            .readdatavalid
		.avm_m1_address       (uart_fast_0_m1_address),                     //            .address
		.avm_m1_writedata     (uart_fast_0_m1_writedata),                   //            .writedata
		.avm_m1_readdata      (uart_fast_0_m1_readdata),                    //            .readdata
		.uart_rx              (uart_rx),                                    // conduit_end.rx
		.uart_tx              (uart_tx)                                     //            .tx
	);

	mySystem_mm_interconnect_0 mm_interconnect_0 (
		.Clock_clk_clk                            (clk_clk),                                                    //                       Clock_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                             // CPU_reset_reset_bridge_in_reset.reset
		.Conclover_0_m1_address                   (conclover_0_m1_address),                                     //                  Conclover_0_m1.address
		.Conclover_0_m1_waitrequest               (conclover_0_m1_waitrequest),                                 //                                .waitrequest
		.Conclover_0_m1_read                      (conclover_0_m1_read),                                        //                                .read
		.Conclover_0_m1_readdata                  (conclover_0_m1_readdata),                                    //                                .readdata
		.Conclover_0_m1_readdatavalid             (conclover_0_m1_readdatavalid),                               //                                .readdatavalid
		.Conclover_0_m1_write                     (conclover_0_m1_write),                                       //                                .write
		.Conclover_0_m1_writedata                 (conclover_0_m1_writedata),                                   //                                .writedata
		.CPU_data_master_address                  (cpu_data_master_address),                                    //                 CPU_data_master.address
		.CPU_data_master_waitrequest              (cpu_data_master_waitrequest),                                //                                .waitrequest
		.CPU_data_master_byteenable               (cpu_data_master_byteenable),                                 //                                .byteenable
		.CPU_data_master_read                     (cpu_data_master_read),                                       //                                .read
		.CPU_data_master_readdata                 (cpu_data_master_readdata),                                   //                                .readdata
		.CPU_data_master_write                    (cpu_data_master_write),                                      //                                .write
		.CPU_data_master_writedata                (cpu_data_master_writedata),                                  //                                .writedata
		.CPU_data_master_debugaccess              (cpu_data_master_debugaccess),                                //                                .debugaccess
		.CPU_instruction_master_address           (cpu_instruction_master_address),                             //          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest       (cpu_instruction_master_waitrequest),                         //                                .waitrequest
		.CPU_instruction_master_read              (cpu_instruction_master_read),                                //                                .read
		.CPU_instruction_master_readdata          (cpu_instruction_master_readdata),                            //                                .readdata
		.UART_Fast_0_m1_address                   (uart_fast_0_m1_address),                                     //                  UART_Fast_0_m1.address
		.UART_Fast_0_m1_waitrequest               (uart_fast_0_m1_waitrequest),                                 //                                .waitrequest
		.UART_Fast_0_m1_read                      (uart_fast_0_m1_read),                                        //                                .read
		.UART_Fast_0_m1_readdata                  (uart_fast_0_m1_readdata),                                    //                                .readdata
		.UART_Fast_0_m1_readdatavalid             (uart_fast_0_m1_readdatavalid),                               //                                .readdatavalid
		.UART_Fast_0_m1_write                     (uart_fast_0_m1_write),                                       //                                .write
		.UART_Fast_0_m1_writedata                 (uart_fast_0_m1_writedata),                                   //                                .writedata
		.Conclover_0_s0_address                   (mm_interconnect_0_conclover_0_s0_address),                   //                  Conclover_0_s0.address
		.Conclover_0_s0_write                     (mm_interconnect_0_conclover_0_s0_write),                     //                                .write
		.Conclover_0_s0_read                      (mm_interconnect_0_conclover_0_s0_read),                      //                                .read
		.Conclover_0_s0_readdata                  (mm_interconnect_0_conclover_0_s0_readdata),                  //                                .readdata
		.Conclover_0_s0_writedata                 (mm_interconnect_0_conclover_0_s0_writedata),                 //                                .writedata
		.CPU_debug_mem_slave_address              (mm_interconnect_0_cpu_debug_mem_slave_address),              //             CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write                (mm_interconnect_0_cpu_debug_mem_slave_write),                //                                .write
		.CPU_debug_mem_slave_read                 (mm_interconnect_0_cpu_debug_mem_slave_read),                 //                                .read
		.CPU_debug_mem_slave_readdata             (mm_interconnect_0_cpu_debug_mem_slave_readdata),             //                                .readdata
		.CPU_debug_mem_slave_writedata            (mm_interconnect_0_cpu_debug_mem_slave_writedata),            //                                .writedata
		.CPU_debug_mem_slave_byteenable           (mm_interconnect_0_cpu_debug_mem_slave_byteenable),           //                                .byteenable
		.CPU_debug_mem_slave_waitrequest          (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),          //                                .waitrequest
		.CPU_debug_mem_slave_debugaccess          (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),          //                                .debugaccess
		.Debug_UART_avalon_jtag_slave_address     (mm_interconnect_0_debug_uart_avalon_jtag_slave_address),     //    Debug_UART_avalon_jtag_slave.address
		.Debug_UART_avalon_jtag_slave_write       (mm_interconnect_0_debug_uart_avalon_jtag_slave_write),       //                                .write
		.Debug_UART_avalon_jtag_slave_read        (mm_interconnect_0_debug_uart_avalon_jtag_slave_read),        //                                .read
		.Debug_UART_avalon_jtag_slave_readdata    (mm_interconnect_0_debug_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.Debug_UART_avalon_jtag_slave_writedata   (mm_interconnect_0_debug_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.Debug_UART_avalon_jtag_slave_waitrequest (mm_interconnect_0_debug_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.Debug_UART_avalon_jtag_slave_chipselect  (mm_interconnect_0_debug_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.Input_s0_address                         (mm_interconnect_0_input_s0_address),                         //                        Input_s0.address
		.Input_s0_write                           (mm_interconnect_0_input_s0_write),                           //                                .write
		.Input_s0_read                            (mm_interconnect_0_input_s0_read),                            //                                .read
		.Input_s0_readdata                        (mm_interconnect_0_input_s0_readdata),                        //                                .readdata
		.Input_s0_writedata                       (mm_interconnect_0_input_s0_writedata),                       //                                .writedata
		.RAM_s1_address                           (mm_interconnect_0_ram_s1_address),                           //                          RAM_s1.address
		.RAM_s1_write                             (mm_interconnect_0_ram_s1_write),                             //                                .write
		.RAM_s1_readdata                          (mm_interconnect_0_ram_s1_readdata),                          //                                .readdata
		.RAM_s1_writedata                         (mm_interconnect_0_ram_s1_writedata),                         //                                .writedata
		.RAM_s1_byteenable                        (mm_interconnect_0_ram_s1_byteenable),                        //                                .byteenable
		.RAM_s1_chipselect                        (mm_interconnect_0_ram_s1_chipselect),                        //                                .chipselect
		.RAM_s1_clken                             (mm_interconnect_0_ram_s1_clken),                             //                                .clken
		.Seven_Segment_Display_s0_address         (mm_interconnect_0_seven_segment_display_s0_address),         //        Seven_Segment_Display_s0.address
		.Seven_Segment_Display_s0_write           (mm_interconnect_0_seven_segment_display_s0_write),           //                                .write
		.Seven_Segment_Display_s0_read            (mm_interconnect_0_seven_segment_display_s0_read),            //                                .read
		.Seven_Segment_Display_s0_readdata        (mm_interconnect_0_seven_segment_display_s0_readdata),        //                                .readdata
		.Seven_Segment_Display_s0_writedata       (mm_interconnect_0_seven_segment_display_s0_writedata),       //                                .writedata
		.System_Timer_s0_address                  (mm_interconnect_0_system_timer_s0_address),                  //                 System_Timer_s0.address
		.System_Timer_s0_write                    (mm_interconnect_0_system_timer_s0_write),                    //                                .write
		.System_Timer_s0_read                     (mm_interconnect_0_system_timer_s0_read),                     //                                .read
		.System_Timer_s0_readdata                 (mm_interconnect_0_system_timer_s0_readdata),                 //                                .readdata
		.System_Timer_s0_writedata                (mm_interconnect_0_system_timer_s0_writedata),                //                                .writedata
		.UART_Fast_0_s0_address                   (mm_interconnect_0_uart_fast_0_s0_address),                   //                  UART_Fast_0_s0.address
		.UART_Fast_0_s0_write                     (mm_interconnect_0_uart_fast_0_s0_write),                     //                                .write
		.UART_Fast_0_s0_read                      (mm_interconnect_0_uart_fast_0_s0_read),                      //                                .read
		.UART_Fast_0_s0_readdata                  (mm_interconnect_0_uart_fast_0_s0_readdata),                  //                                .readdata
		.UART_Fast_0_s0_writedata                 (mm_interconnect_0_uart_fast_0_s0_writedata)                  //                                .writedata
	);

	mySystem_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
